.subckt ecg n1 n2				
vin n1 n2 pwl				
+	0.0001	0.84934663		
+	0.0002	0.86012948		
+	0.0003	0.88099758		
+	0.0004	0.88138071		
+	0.0005	0.8782381		
+	0.0006	0.87514976		
+	0.0007	0.88580609		
+	0.0008	0.88444072		
+	0.0009	0.89321629		
+	0.001	0.88178824		
+	0.0011	0.88994316		
+	0.0012	0.88955006		
+	0.0013	0.89383242		
+	0.0014	0.88543983		
+	0.0015	0.88732395		
+	0.0016	0.90098087		
+	0.0017	0.91044309		
+	0.0018	0.89772692		
+	0.0019	0.9105633		
+	0.002	0.91836327		
+	0.0021	0.91400666		
+	0.0022	0.9241377		
+	0.0023	0.9135295		
+	0.0024	0.92643908		
+	0.0025	0.91982628		
+	0.0026	0.91714282		
+	0.0027	0.93814095		
+	0.0028	0.92773108		
+	0.0029	0.94693186		
+	0.003	0.95004493		
+	0.0031	0.96147651		
+	0.0032	0.96913823		
+	0.0033	0.98216212		
+	0.0034	0.97111864		
+	0.0035	0.97402266		
+	0.0036	0.97415236		
+	0.0037	0.96771027		
+	0.0038	0.97456181		
+	0.0039	0.97388006		
+	0.004	0.978335		
+	0.0041	0.96078967		
+	0.0042	0.96018427		
+	0.0043	0.95551332		
+	0.0044	0.96014455		
+	0.0045	0.95616897		
+	0.0046	0.94190751		
+	0.0047	0.93884085		
+	0.0048	0.94341827		
+	0.0049	0.946374		
+	0.005	0.93113991		
+	0.0051	0.93652093		
+	0.0052	0.93498496		
+	0.0053	0.94229587		
+	0.0054	0.92824146		
+	0.0055	0.93182816		
+	0.0056	0.9482858		
+	0.0057	0.94105171		
+	0.0058	0.95150803		
+	0.0059	0.96484336		
+	0.006	0.98301147		
+	0.0061	0.98213388		
+	0.0062	0.99001126		
+	0.0063	0.99488558		
+	0.0064	0.98264383		
+	0.0065	0.98432741		
+	0.0066	0.98680065		
+	0.0067	0.97420028		
+	0.0068	0.97257417		
+	0.0069	0.96846235		
+	0.007	0.97546497		
+	0.0071	0.96333275		
+	0.0072	0.95954651		
+	0.0073	0.94708182		
+	0.0074	0.93778489		
+	0.0075	0.93119208		
+	0.0076	0.90326348		
+	0.0077	0.90722793		
+	0.0078	0.89383384		
+	0.0079	0.87913513		
+	0.008	0.87551099		
+	0.0081	0.8763784		
+	0.0082	0.8672192		
+	0.0083	0.86570546		
+	0.0084	0.84843747		
+	0.0085	0.85498422		
+	0.0086	0.84974363		
+	0.0087	0.85556179		
+	0.0088	0.86496661		
+	0.0089	0.88023365		
+	0.009	0.88473828		
+	0.0091	0.88954507		
+	0.0092	0.88075561		
+	0.0093	0.88602876		
+	0.0094	0.87878353		
+	0.0095	0.87542498		
+	0.0096	0.86534305		
+	0.0097	0.87505189		
+	0.0098	0.86692341		
+	0.0099	0.86263038		
+	0.01	0.85624204		
+	0.0101	0.86203364		
+	0.0102	0.8446523		
+	0.0103	0.84025058		
+	0.0104	0.83281588		
+	0.0105	0.83384531		
+	0.0106	0.84452596		
+	0.0107	0.83129826		
+	0.0108	0.83151202		
+	0.0109	0.82272155		
+	0.011	0.83307705		
+	0.0111	0.81742778		
+	0.0112	0.82035897		
+	0.0113	0.82723979		
+	0.0114	0.81806908		
+	0.0115	0.82995629		
+	0.0116	0.84893364		
+	0.0117	0.85515527		
+	0.0118	0.86390635		
+	0.0119	0.87309616		
+	0.012	0.87470586		
+	0.0121	0.87302748		
+	0.0122	0.88004523		
+	0.0123	0.86763893		
+	0.0124	0.8697488		
+	0.0125	0.8791125		
+	0.0126	0.86440952		
+	0.0127	0.87722939		
+	0.0128	0.86159762		
+	0.0129	0.86332318		
+	0.013	0.85710807		
+	0.0131	0.84861945		
+	0.0132	0.8466127		
+	0.0133	0.85403973		
+	0.0134	0.84803914		
+	0.0135	0.83579578		
+	0.0136	0.84586849		
+	0.0137	0.82571621		
+	0.0138	0.83878578		
+	0.0139	0.83945027		
+	0.014	0.82641209		
+	0.0141	0.82718059		
+	0.0142	0.82061108		
+	0.0143	0.82874075		
+	0.0144	0.82543358		
+	0.0145	0.83598482		
+	0.0146	0.86175669		
+	0.0147	0.86473651		
+	0.0148	0.87175707		
+	0.0149	0.87187262		
+	0.015	0.88199112		
+	0.0151	0.8812959		
+	0.0152	0.87472951		
+	0.0153	0.88371576		
+	0.0154	0.87383907		
+	0.0155	0.877698		
+	0.0156	0.87141423		
+	0.0157	0.86727546		
+	0.0158	0.86306131		
+	0.0159	0.866797		
+	0.016	0.85176573		
+	0.0161	0.85061751		
+	0.0162	0.84621909		
+	0.0163	0.84174703		
+	0.0164	0.84108651		
+	0.0165	0.84277697		
+	0.0166	0.84159888		
+	0.0167	0.84924397		
+	0.0168	0.85128144		
+	0.0169	0.84586731		
+	0.017	0.84650899		
+	0.0171	0.85704503		
+	0.0172	0.84999745		
+	0.0173	0.85433392		
+	0.0174	0.87631409		
+	0.0175	0.88922903		
+	0.0176	0.9029057		
+	0.0177	0.93208343		
+	0.0178	0.94723825		
+	0.0179	0.94891789		
+	0.018	0.949071		
+	0.0181	0.96609913		
+	0.0182	0.97169376		
+	0.0183	0.97501335		
+	0.0184	0.96978961		
+	0.0185	0.97283958		
+	0.0186	0.97455651		
+	0.0187	0.97911257		
+	0.0188	0.97655597		
+	0.0189	0.96494314		
+	0.019	0.95791053		
+	0.0191	0.96662752		
+	0.0192	0.96152946		
+	0.0193	0.94634697		
+	0.0194	0.95586402		
+	0.0195	0.95226973		
+	0.0196	0.93911531		
+	0.0197	0.94811703		
+	0.0198	0.93509726		
+	0.0199	0.9403681		
+	0.02	0.94321358		
+	0.0201	0.93835687		
+	0.0202	0.94061058		
+	0.0203	0.94342754		
+	0.0204	0.96604423		
+	0.0205	0.97638568		
+	0.0206	0.99330916		
+	0.0207	0.99382547		
+	0.0208	1.0019221		
+	0.0209	1.0053997		
+	0.021	0.98751199		
+	0.0211	0.9968252		
+	0.0212	0.99804445		
+	0.0213	0.99779839		
+	0.0214	0.98921192		
+	0.0215	0.98858291		
+	0.0216	0.98772417		
+	0.0217	0.97545437		
+	0.0218	0.98314744		
+	0.0219	0.96466598		
+	0.022	0.96414426		
+	0.0221	0.97290278		
+	0.0222	0.95923536		
+	0.0223	0.95605623		
+	0.0224	0.95638128		
+	0.0225	0.94757521		
+	0.0226	0.94663575		
+	0.0227	0.95887845		
+	0.0228	0.94974322		
+	0.0229	0.94245165		
+	0.023	0.93834069		
+	0.0231	0.94839382		
+	0.0232	0.94926094		
+	0.0233	0.9639264		
+	0.0234	0.96647886		
+	0.0235	0.9779951		
+	0.0236	0.96997086		
+	0.0237	0.9704953		
+	0.0238	0.95447384		
+	0.0239	0.95923362		
+	0.024	0.94036098		
+	0.0241	0.93377722		
+	0.0242	0.93807193		
+	0.0243	0.92112418		
+	0.0244	0.91879834		
+	0.0245	0.91408166		
+	0.0246	0.89972898		
+	0.0247	0.88445927		
+	0.0248	0.87993527		
+	0.0249	0.87128714		
+	0.025	0.86642856		
+	0.0251	0.87143918		
+	0.0252	0.85044367		
+	0.0253	0.86407705		
+	0.0254	0.85775333		
+	0.0255	0.83727454		
+	0.0256	0.83761634		
+	0.0257	0.83319057		
+	0.0258	0.83568139		
+	0.0259	0.82738828		
+	0.026	0.83373496		
+	0.0261	0.84851088		
+	0.0262	0.85789724		
+	0.0263	0.86598384		
+	0.0264	0.86748123		
+	0.0265	0.87412555		
+	0.0266	0.88676978		
+	0.0267	0.87976495		
+	0.0268	0.89062735		
+	0.0269	0.88344032		
+	0.027	0.89221423		
+	0.0271	0.88097276		
+	0.0272	0.87264977		
+	0.0273	0.86777569		
+	0.0274	0.86536591		
+	0.0275	0.86581193		
+	0.0276	0.86396089		
+	0.0277	0.8651437		
+	0.0278	0.85523856		
+	0.0279	0.86444145		
+	0.028	0.84459212		
+	0.0281	0.84933133		
+	0.0282	0.84573436		
+	0.0283	0.85034487		
+	0.0284	0.84953874		
+	0.0285	0.84845044		
+	0.0286	0.83324994		
+	0.0287	0.84111458		
+	0.0288	0.83518942		
+	0.0289	0.83591577		
+	0.029	0.85047379		
+	0.0291	0.85739362		
+	0.0292	0.85577884		
+	0.0293	0.86505607		
+	0.0294	0.86876868		
+	0.0295	0.8893719		
+	0.0296	0.87878162		
+	0.0297	0.89773904		
+	0.0298	0.88145516		
+	0.0299	0.89566517		
+	0.03	0.8903824		
+	0.0301	0.88362579		
+	0.0302	0.88390253		
+	0.0303	0.87617527		
+	0.0304	0.86663823		
+	0.0305	0.86250666		
+	0.0306	0.86517256		
+	0.0307	0.87130895		
+	0.0308	0.85743425		
+	0.0309	0.86347381		
+	0.031	0.85599524		
+	0.0311	0.85482153		
+	0.0312	0.84437877		
+	0.0313	0.8536997		
+	0.0314	0.85013239		
+	0.0315	0.84852744		
+	0.0316	0.84397191		
+	0.0317	0.83412133		
+	0.0318	0.84282462		
+	0.0319	0.83483236		
+	0.032	0.8395685		
+	0.0321	0.86861606		
+	0.0322	0.87571503		
+	0.0323	0.88777517		
+	0.0324	0.88446732		
+	0.0325	0.88662863		
+	0.0326	0.89919086		
+	0.0327	0.89125695		
+	0.0328	0.89375417		
+	0.0329	0.89059183		
+	0.033	0.88864818		
+	0.0331	0.88615144		
+	0.0332	0.89544216		
+	0.0333	0.9058001		
+	0.0334	0.90695709		
+	0.0335	0.90481389		
+	0.0336	0.89898778		
+	0.0337	0.90844183		
+	0.0338	0.91484694		
+	0.0339	0.91281233		
+	0.034	0.90827537		
+	0.0341	0.9117027		
+	0.0342	0.90935939		
+	0.0343	0.92213464		
+	0.0344	0.92279916		
+	0.0345	0.9250502		
+	0.0346	0.92707024		
+	0.0347	0.94637156		
+	0.0348	0.94314874		
+	0.0349	0.94491626		
+	0.035	0.95981782		
+	0.0351	0.96784998		
+	0.0352	0.97761662		
+	0.0353	0.99478998		
+	0.0354	0.99647092		
+	0.0355	0.99321086		
+	0.0356	0.98921662		
+	0.0357	0.98907638		
+	0.0358	0.99759239		
+	0.0359	0.98807394		
+	0.036	0.9932705		
+	0.0361	0.9945637		
+	0.0362	0.9984927		
+	0.0363	0.98746497		
+	0.0364	0.98737771		
+	0.0365	0.98387083		
+	0.0366	0.97325019		
+	0.0367	0.9741259		
+	0.0368	0.9715199		
+	0.0369	0.97525512		
+	0.037	0.97352078		
+	0.0371	0.96912767		
+	0.0372	0.95310406		
+	0.0373	0.95490403		
+	0.0374	0.95750552		
+	0.0375	0.96066631		
+	0.0376	0.95050263		
+	0.0377	0.96301603		
+	0.0378	0.96600847		
+	0.0379	0.97013927		
+	0.038	0.97410796		
+	0.0381	0.98762474		
+	0.0382	0.99774006		
+	0.0383	1.0008392		
+	0.0384	1.0116725		
+	0.0385	1.0114857		
+	0.0386	1.0106765		
+	0.0387	1.0016319		
+	0.0388	1.0131608		
+	0.0389	1.0013278		
+	0.039	1.0034544		
+	0.0391	1.0000679		
+	0.0392	0.99583047		
+	0.0393	0.98150545		
+	0.0394	0.98283294		
+	0.0395	0.98227363		
+	0.0396	0.9638498		
+	0.0397	0.97001127		
+	0.0398	0.95771838		
+	0.0399	0.93892463		
+	0.04	0.93624586		
+	0.0401	0.92245278		
+	0.0402	0.91291488		
+	0.0403	0.89279018		
+	0.0404	0.90206616		
+	0.0405	0.8804997		
+	0.0406	0.8924684		
+	0.0407	0.89215217		
+	0.0408	0.88603464		
+	0.0409	0.89239133		
+	0.041	0.90478176		
+	0.0411	0.90739508		
+	0.0412	0.91584749		
+	0.0413	0.91030863		
+	0.0414	0.90153465		
+	0.0415	0.90077516		
+	0.0416	0.90753539		
+	0.0417	0.90700161		
+	0.0418	0.88577482		
+	0.0419	0.88091063		
+	0.042	0.88042378		
+	0.0421	0.87404131		
+	0.0422	0.88145111		
+	0.0423	0.86733574		
+	0.0424	0.87799498		
+	0.0425	0.85574019		
+	0.0426	0.85753504		
+	0.0427	0.85389553		
+	0.0428	0.84577533		
+	0.0429	0.8602717		
+	0.043	0.84665335		
+	0.0431	0.85486096		
+	0.0432	0.84575567		
+	0.0433	0.8494496		
+	0.0434	0.83567907		
+	0.0435	0.8472366		
+	0.0436	0.83787398		
+	0.0437	0.84752245		
+	0.0438	0.85833396		
+	0.0439	0.88239356		
+	0.044	0.89010943		
+	0.0441	0.88570275		
+	0.0442	0.89363783		
+	0.0443	0.89864035		
+	0.0444	0.89953936		
+	0.0445	0.89649614		
+	0.0446	0.89088938		
+	0.0447	0.88605953		
+	0.0448	0.89074869		
+	0.0449	0.87935828		
+	0.045	0.88677134		
+	0.0451	0.88287674		
+	0.0452	0.86760391		
+	0.0453	0.87937887		
+	0.0454	0.86580677		
+	0.0455	0.85750709		
+	0.0456	0.86170026		
+	0.0457	0.86664705		
+	0.0458	0.85328663		
+	0.0459	0.85713107		
+	0.046	0.84867396		
+	0.0461	0.85161621		
+	0.0462	0.84095454		
+	0.0463	0.84054		
+	0.0464	0.85518753		
+	0.0465	0.85482642		
+	0.0466	0.84925976		
+	0.0467	0.86871677		
+	0.0468	0.87468586		
+	0.0469	0.88159021		
+	0.047	0.90010695		
+	0.0471	0.89350623		
+	0.0472	0.90019772		
+	0.0473	0.89783905		
+	0.0474	0.90530542		
+	0.0475	0.88674804		
+	0.0476	0.89648487		
+	0.0477	0.89259335		
+	0.0478	0.89398923		
+	0.0479	0.88426247		
+	0.048	0.88274229		
+	0.0481	0.8860524		
+	0.0482	0.88210167		
+	0.0483	0.86810127		
+	0.0484	0.86072142		
+	0.0485	0.86002741		
+	0.0486	0.8599625		
+	0.0487	0.85022577		
+	0.0488	0.85400814		
+	0.0489	0.85932734		
+	0.049	0.85635325		
+	0.0491	0.86331591		
+	0.0492	0.85241827		
+	0.0493	0.86490519		
+	0.0494	0.86043835		
+	0.0495	0.8697959		
+	0.0496	0.88546624		
+	0.0497	0.89929338		
+	0.0498	0.90901473		
+	0.0499	0.94140256		
+	0.05	0.94896813		
+	0.0501	0.94539353		
+	0.0502	0.95719904		
+	0.0503	0.96931694		
+	0.0504	0.96076454		
+	0.0505	0.970512		
+	0.0506	0.97861704		
+	0.0507	0.97204953		
+	0.0508	0.98112572		
+	0.0509	0.98358458		
+	0.051	0.97007322		
+	0.0511	0.98230267		
+	0.0512	0.97854845		
+	0.0513	0.98012541		
+	0.0514	0.96351927		
+	0.0515	0.96760053		
+	0.0516	0.9695151		
+	0.0517	0.958758		
+	0.0518	0.95178299		
+	0.0519	0.95523035		
+	0.052	0.96747238		
+	0.0521	0.94998704		
+	0.0522	0.95585092		
+	0.0523	0.96425837		
+	0.0524	0.96248517		
+	0.0525	0.97308233		
+	0.0526	0.98764051		
+	0.0527	0.98497047		
+	0.0528	0.99459591		
+	0.0529	1.0186421		
+	0.053	1.0208472		
+	0.0531	1.0036277		
+	0.0532	1.0210984		
+	0.0533	1.0189623		
+	0.0534	1.014336		
+	0.0535	1.0132938		
+	0.0536	1.0024625		
+	0.0537	0.99851525		
+	0.0538	0.99843083		
+	0.0539	1.0018013		
+	0.054	0.99583962		
+	0.0541	0.98834473		
+	0.0542	0.98913265		
+	0.0543	0.97576677		
+	0.0544	0.9823955		
+	0.0545	0.97749563		
+	0.0546	0.96678029		
+	0.0547	0.96093499		
+	0.0548	0.96989924		
+	0.0549	0.96212648		
+	0.055	0.96778923		
+	0.0551	0.95838031		
+	0.0552	0.96887818		
+	0.0553	0.96365622		
+	0.0554	0.9683736		
+	0.0555	0.97987347		
+	0.0556	0.99680839		
+	0.0557	1.0043219		
+	0.0558	0.99345638		
+	0.0559	1.0026573		
+	0.056	0.99981695		
+	0.0561	0.98907052		
+	0.0562	0.97343035		
+	0.0563	0.961964		
+	0.0564	0.96214182		
+	0.0565	0.95589001		
+	0.0566	0.93815946		
+	0.0567	0.93040705		
+	0.0568	0.92156989		
+	0.0569	0.92095395		
+	0.057	0.91213169		
+	0.0571	0.90152705		
+	0.0572	0.89537255		
+	0.0573	0.89447574		
+	0.0574	0.8805148		
+	0.0575	0.88432625		
+	0.0576	0.87007251		
+	0.0577	0.86398778		
+	0.0578	0.86638719		
+	0.0579	0.84839792		
+	0.058	0.85126403		
+	0.0581	0.85734625		
+	0.0582	0.86492657		
+	0.0583	0.85883658		
+	0.0584	0.87442962		
+	0.0585	0.88374686		
+	0.0586	0.89701257		
+	0.0587	0.89742157		
+	0.0588	0.90783867		
+	0.0589	0.89567919		
+	0.059	0.9072055		
+	0.0591	0.8941315		
+	0.0592	0.89811848		
+	0.0593	0.90401729		
+	0.0594	0.90206463		
+	0.0595	0.89926399		
+	0.0596	0.88634239		
+	0.0597	0.88477779		
+	0.0598	0.88243045		
+	0.0599	0.88371948		
+	0.06	0.87007933		
+	0.0601	0.87531766		
+	0.0602	0.87136421		
+	0.0603	0.86083221		
+	0.0604	0.85847956		
+	0.0605	0.86341126		
+	0.0606	0.85855655		
+	0.0607	0.85159764		
+	0.0608	0.84900577		
+	0.0609	0.84199899		
+	0.061	0.84405669		
+	0.0611	0.85485113		
+	0.0612	0.85466853		
+	0.0613	0.85885236		
+	0.0614	0.87667862		
+	0.0615	0.88359468		
+	0.0616	0.88876218		
+	0.0617	0.90108866		
+	0.0618	0.89337983		
+	0.0619	0.90309782		
+	0.062	0.90120632		
+	0.0621	0.89934796		
+	0.0622	0.89507119		
+	0.0623	0.89047944		
+	0.0624	0.89505841		
+	0.0625	0.88574865		
+	0.0626	0.88425565		
+	0.0627	0.8857759		
+	0.0628	0.878188		
+	0.0629	0.87042111		
+	0.063	0.88129077		
+	0.0631	0.8648184		
+	0.0632	0.86019662		
+	0.0633	0.85774451		
+	0.0634	0.85013983		
+	0.0635	0.85628184		
+	0.0636	0.865366		
+	0.0637	0.85733669		
+	0.0638	0.84808185		
+	0.0639	0.85190178		
+	0.064	0.84766824		
+	0.0641	0.85256883		
+	0.0642	0.87351457		
+	0.0643	0.88151758		
+	0.0644	0.87743068		
+	0.0645	0.89367675		
+	0.0646	0.90221935		
+	0.0647	0.91274856		
+	0.0648	0.91046466		
+	0.0649	0.91097152		
+	0.065	0.90717258		
+	0.0651	0.90933916		
+	0.0652	0.91229334		
+	0.0653	0.89301002		
+	0.0654	0.89588069		
+	0.0655	0.89697885		
+	0.0656	0.90460743		
+	0.0657	0.90179915		
+	0.0658	0.89779701		
+	0.0659	0.9083126		
+	0.066	0.90296983		
+	0.0661	0.90605288		
+	0.0662	0.91764609		
+	0.0663	0.90784293		
+	0.0664	0.9091655		
+	0.0665	0.91330976		
+	0.0666	0.92444872		
+	0.0667	0.93225042		
+	0.0668	0.94406514		
+	0.0669	0.93199227		
+	0.067	0.95023788		
+	0.0671	0.96327911		
+	0.0672	0.96594452		
+	0.0673	0.99068467		
+	0.0674	0.98640893		
+	0.0675	0.99929117		
+	0.0676	1.0093096		
+	0.0677	1.0138648		
+	0.0678	1.0145851		
+	0.0679	1.0043296		
+	0.068	1.0063478		
+	0.0681	1.0130399		
+	0.0682	1.0008691		
+	0.0683	0.99351492		
+	0.0684	0.99045172		
+	0.0685	0.9912022		
+	0.0686	0.9941811		
+	0.0687	0.99508592		
+	0.0688	0.98379928		
+	0.0689	0.98717157		
+	0.069	0.98597589		
+	0.0691	0.97801338		
+	0.0692	0.97484378		
+	0.0693	0.97233185		
+	0.0694	0.96369148		
+	0.0695	0.9629179		
+	0.0696	0.96649629		
+	0.0697	0.96377555		
+	0.0698	0.97116529		
+	0.0699	0.97435498		
+	0.07	0.98414391		
+	0.0701	0.97779231		
+	0.0702	0.99921287		
+	0.0703	1.007552		
+	0.0704	1.0181981		
+	0.0705	1.0257221		
+	0.0706	1.0276318		
+	0.0707	1.0265525		
+	0.0708	1.0218011		
+	0.0709	1.022797		
+	0.071	1.0101189		
+	0.0711	1.0055337		
+	0.0712	1.0072645		
+	0.0713	0.99772686		
+	0.0714	1.0030011		
+	0.0715	1.0049476		
+	0.0716	0.99006171		
+	0.0717	0.98686674		
+	0.0718	0.9913741		
+	0.0719	0.98178419		
+	0.072	0.97556435		
+	0.0721	0.97279932		
+	0.0722	0.95152071		
+	0.0723	0.95208761		
+	0.0724	0.94134052		
+	0.0725	0.93641329		
+	0.0726	0.91791504		
+	0.0727	0.9110313		
+	0.0728	0.91446733		
+	0.0729	0.9032002		
+	0.073	0.90654783		
+	0.0731	0.91398154		
+	0.0732	0.91500469		
+	0.0733	0.93570204		
+	0.0734	0.92306762		
+	0.0735	0.92861483		
+	0.0736	0.92839988		
+	0.0737	0.91690647		
+	0.0738	0.91056934		
+	0.0739	0.91091946		
+	0.074	0.89920644		
+	0.0741	0.90596982		
+	0.0742	0.90852205		
+	0.0743	0.89529231		
+	0.0744	0.89631938		
+	0.0745	0.88012431		
+	0.0746	0.87845952		
+	0.0747	0.86894235		
+	0.0748	0.86046736		
+	0.0749	0.87426986		
+	0.075	0.86820691		
+	0.0751	0.85707761		
+	0.0752	0.8623189		
+	0.0753	0.84937607		
+	0.0754	0.84559523		
+	0.0755	0.85540763		
+	0.0756	0.85816647		
+	0.0757	0.85388244		
+	0.0758	0.85689876		
+	0.0759	0.87586291		
+	0.076	0.87211336		
+	0.0761	0.89283971		
+	0.0762	0.90068961		
+	0.0763	0.89724182		
+	0.0764	0.90055136		
+	0.0765	0.91008128		
+	0.0766	0.90589916		
+	0.0767	0.91166754		
+	0.0768	0.89428423		
+	0.0769	0.89457463		
+	0.077	0.89513329		
+	0.0771	0.8871196		
+	0.0772	0.89756769		
+	0.0773	0.88896732		
+	0.0774	0.8880343		
+	0.0775	0.88083801		
+	0.0776	0.86608062		
+	0.0777	0.87925943		
+	0.0778	0.87637191		
+	0.0779	0.85968032		
+	0.078	0.86816159		
+	0.0781	0.8568773		
+	0.0782	0.85503468		
+	0.0783	0.85921278		
+	0.0784	0.84931616		
+	0.0785	0.85733932		
+	0.0786	0.85900911		
+	0.0787	0.86485692		
+	0.0788	0.8702034		
+	0.0789	0.87528716		
+	0.079	0.87636709		
+	0.0791	0.88863483		
+	0.0792	0.89758491		
+	0.0793	0.90130491		
+	0.0794	0.89964129		
+	0.0795	0.90600097		
+	0.0796	0.89609155		
+	0.0797	0.89358971		
+	0.0798	0.90792473		
+	0.0799	0.89119763		
+	0.08	0.89382087		
+	0.0801	0.89213271		
+	0.0802	0.88574332		
+	0.0803	0.88546941		
+	0.0804	0.87725278		
+	0.0805	0.88365472		
+	0.0806	0.86694514		
+	0.0807	0.86828721		
+	0.0808	0.86206242		
+	0.0809	0.87379817		
+	0.081	0.86223968		
+	0.0811	0.86063692		
+	0.0812	0.86540704		
+	0.0813	0.84982109		
+	0.0814	0.85257374		
+	0.0815	0.86450974		
+	0.0816	0.85878725		
+	0.0817	0.86821421		
+	0.0818	0.8862221		
+	0.0819	0.90687577		
+	0.082	0.91560174		
+	0.0821	0.91972677		
+	0.0822	0.93292984		
+	0.0823	0.95306043		
+	0.0824	0.94866464		
+	0.0825	0.95853809		
+	0.0826	0.96157056		
+	0.0827	0.96763367		
+	0.0828	0.96896564		
+	0.0829	0.9761487		
+	0.083	0.98469324		
+	0.0831	0.98429464		
+	0.0832	0.97165807		
+	0.0833	0.97976494		
+	0.0834	0.96938756		
+	0.0835	0.97156616		
+	0.0836	0.97203242		
+	0.0837	0.97574135		
+	0.0838	0.96735775		
+	0.0839	0.96726321		
+	0.084	0.96306346		
+	0.0841	0.96738996		
+	0.0842	0.95389866		
+	0.0843	0.9605485		
+	0.0844	0.95687695		
+	0.0845	0.95562367		
+	0.0846	0.9623826		
+	0.0847	0.98420391		
+	0.0848	0.98733898		
+	0.0849	1.0055411		
+	0.085	1.0172531		
+	0.0851	1.0259179		
+	0.0852	1.0192947		
+	0.0853	1.0200178		
+	0.0854	1.0088431		
+	0.0855	1.0243635		
+	0.0856	1.0205508		
+	0.0857	1.0152549		
+	0.0858	1.0079297		
+	0.0859	1.0060767		
+	0.086	1.0033098		
+	0.0861	0.99876279		
+	0.0862	0.99822766		
+	0.0863	0.98638703		
+	0.0864	0.99475366		
+	0.0865	0.98495053		
+	0.0866	0.97976277		
+	0.0867	0.96884626		
+	0.0868	0.98316783		
+	0.0869	0.97477195		
+	0.087	0.96666806		
+	0.0871	0.97518878		
+	0.0872	0.95926147		
+	0.0873	0.97404641		
+	0.0874	0.97494005		
+	0.0875	0.97680683		
+	0.0876	0.9769263		
+	0.0877	0.98566843		
+	0.0878	0.99328871		
+	0.0879	1.0130787		
+	0.088	1.0072997		
+	0.0881	1.0228112		
+	0.0882	1.0113443		
+	0.0883	1.0104145		
+	0.0884	1.0098691		
+	0.0885	1.0015129		
+	0.0886	0.98117251		
+	0.0887	0.97560043		
+	0.0888	0.96600029		
+	0.0889	0.9463747		
+	0.089	0.93469252		
+	0.0891	0.93082917		
+	0.0892	0.91853146		
+	0.0893	0.91606117		
+	0.0894	0.91411733		
+	0.0895	0.90887346		
+	0.0896	0.89019157		
+	0.0897	0.88363761		
+	0.0898	0.88916775		
+	0.0899	0.86751205		
+	0.09	0.8697999		
+	0.0901	0.86823871		
+	0.0902	0.86444304		
+	0.0903	0.85275733		
+	0.0904	0.86425804		
+	0.0905	0.87384529		
+	0.0906	0.87329329		
+	0.0907	0.88908901		
+	0.0908	0.89127483		
+	0.0909	0.90665238		
+	0.091	0.90770583		
+	0.0911	0.89810294		
+	0.0912	0.9048149		
+	0.0913	0.90651438		
+	0.0914	0.9087347		
+	0.0915	0.90310667		
+	0.0916	0.88923098		
+	0.0917	0.89703225		
+	0.0918	0.89485623		
+	0.0919	0.87833418		
+	0.092	0.88490356		
+	0.0921	0.88729179		
+	0.0922	0.87222706		
+	0.0923	0.86342138		
+	0.0924	0.86459139		
+	0.0925	0.87207615		
+	0.0926	0.86437036		
+	0.0927	0.85369888		
+	0.0928	0.86199775		
+	0.0929	0.85533742		
+	0.093	0.85785401		
+	0.0931	0.85393508		
+	0.0932	0.86207847		
+	0.0933	0.84733574		
+	0.0934	0.86432118		
+	0.0935	0.87361139		
+	0.0936	0.89028853		
+	0.0937	0.88699175		
+	0.0938	0.8930137		
+	0.0939	0.90317962		
+	0.094	0.90766829		
+	0.0941	0.9020673		
+	0.0942	0.91250005		
+	0.0943	0.90941613		
+	0.0944	0.8972434		
+	0.0945	0.89671664		
+	0.0946	0.89346316		
+	0.0947	0.89311999		
+	0.0948	0.88190091		
+	0.0949	0.88982765		
+	0.095	0.87688524		
+	0.0951	0.8783532		
+	0.0952	0.87467319		
+	0.0953	0.86356158		
+	0.0954	0.8625881		
+	0.0955	0.87193933		
+	0.0956	0.8604962		
+	0.0957	0.86516175		
+	0.0958	0.85455146		
+	0.0959	0.8567251		
+	0.096	0.84465907		
+	0.0961	0.85807866		
+	0.0962	0.85083489		
+	0.0963	0.86058972		
+	0.0964	0.86417927		
+	0.0965	0.87347914		
+	0.0966	0.90005185		
+	0.0967	0.89369754		
+	0.0968	0.91399867		
+	0.0969	0.91569751		
+	0.097	0.91410307		
+	0.0971	0.89803595		
+	0.0972	0.89531413		
+	0.0973	0.9110507		
+	0.0974	0.89351691		
+	0.0975	0.89627684		
+	0.0976	0.90479412		
+	0.0977	0.88969361		
+	0.0978	0.90075931		
+	0.0979	0.88622929		
+	0.098	0.88952262		
+	0.0981	0.89600138		
+	0.0982	0.88245525		
+	0.0983	0.89551014		
+	0.0984	0.88602286		
+	0.0985	0.88668123		
+	0.0986	0.90278761		
+	0.0987	0.89533144		
+	0.0988	0.91732237		
+	0.0989	0.90904215		
+	0.099	0.92367918		
+	0.0991	0.91930466		
+	0.0992	0.93300294		
+	0.0993	0.95289028		
+	0.0994	0.97525479		
+	0.0995	0.98353346		
+	0.0996	0.98431153		
+	0.0997	1.0045631		
+	0.0998	1.0056546		
+	0.0999	1.0006985		
+	0.1	0.9978889		
+	0.1001	1.0034096		
+	0.1002	1.0088153		
+	0.1003	1.0002755		
+	0.1004	0.99593999		
+	0.1005	0.99217466		
+	0.1006	0.99331044		
+	0.1007	1.0015456		
+	0.1008	0.98778337		
+	0.1009	0.99365087		
+	0.101	0.98405929		
+	0.1011	0.97962224		
+	0.1012	0.9746012		
+	0.1013	0.98233417		
+	0.1014	0.97951615		
+	0.1015	0.97604611		
+	0.1016	0.97764474		
+	0.1017	0.95771967		
+	0.1018	0.96996793		
+	0.1019	0.97444609		
+	0.102	0.96233684		
+	0.1021	0.97616288		
+	0.1022	0.98476555		
+	0.1023	0.99090532		
+	0.1024	1.0003628		
+	0.1025	1.0099517		
+	0.1026	1.0052981		
+	0.1027	1.0121433		
+	0.1028	1.0248498		
+	0.1029	1.0117122		
+	0.103	1.0064586		
+	0.1031	1.0225348		
+	0.1032	1.0081365		
+	0.1033	1.0135612		
+	0.1034	1.0130296		
+	0.1035	1.0036642		
+	0.1036	1.0055253		
+	0.1037	0.99128157		
+	0.1038	0.98772893		
+	0.1039	0.99060345		
+	0.104	0.97719887		
+	0.1041	0.97005986		
+	0.1042	0.98287291		
+	0.1043	0.96520014		
+	0.1044	0.9667874		
+	0.1045	0.96925897		
+	0.1046	0.95524996		
+	0.1047	0.95165816		
+	0.1048	0.93255654		
+	0.1049	0.9360509		
+	0.105	0.91705683		
+	0.1051	0.91891802		
+	0.1052	0.93576976		
+	0.1053	0.93828743		
+	0.1054	0.94130003		
+	0.1055	0.94982098		
+	0.1056	0.94710383		
+	0.1057	0.93967815		
+	0.1058	0.92828614		
+	0.1059	0.93379838		
+	0.106	0.92325617		
+	0.1061	0.92026093		
+	0.1062	0.90233272		
+	0.1063	0.91538681		
+	0.1064	0.907913		
+	0.1065	0.89155014		
+	0.1066	0.8964705		
+	0.1067	0.88170936		
+	0.1068	0.87305272		
+	0.1069	0.86851124		
+	0.107	0.87305102		
+	0.1071	0.8574815		
+	0.1072	0.86410003		
+	0.1073	0.8590001		
+	0.1074	0.85968922		
+	0.1075	0.84978193		
+	0.1076	0.84257796		
+	0.1077	0.84196599		
+	0.1078	0.8512177		
+	0.1079	0.85734684		
+	0.108	0.84839482		
+	0.1081	0.86327106		
+	0.1082	0.88508141		
+	0.1083	0.88498108		
+	0.1084	0.89883249		
+	0.1085	0.89830762		
+	0.1086	0.90610668		
+	0.1087	0.89769164		
+	0.1088	0.89309321		
+	0.1089	0.90104134		
+	0.109	0.89136463		
+	0.1091	0.89502741		
+	0.1092	0.89566808		
+	0.1093	0.88489887		
+	0.1094	0.87600025		
+	0.1095	0.88372021		
+	0.1096	0.87617228		
+	0.1097	0.87717788		
+	0.1098	0.87311168		
+	0.1099	0.86954655		
+	0.11	0.85722309		
+	0.1101	0.86822097		
+	0.1102	0.84942142		
+	0.1103	0.8485135		
+	0.1104	0.84445973		
+	0.1105	0.84303547		
+	0.1106	0.85096447		
+	0.1107	0.85189584		
+	0.1108	0.85825264		
+	0.1109	0.85742277		
+	0.111	0.86485456		
+	0.1111	0.86905523		
+	0.1112	0.88576001		
+	0.1113	0.90046725		
+	0.1114	0.90426184		
+	0.1115	0.9077307		
+	0.1116	0.91039486		
+	0.1117	0.90654961		
+	0.1118	0.90613009		
+	0.1119	0.90623753		
+	0.112	0.89441633		
+	0.1121	0.88916881		
+	0.1122	0.89786219		
+	0.1123	0.88298051		
+	0.1124	0.8777355		
+	0.1125	0.87616784		
+	0.1126	0.88272937		
+	0.1127	0.86441216		
+	0.1128	0.86043697		
+	0.1129	0.86631815		
+	0.113	0.86997994		
+	0.1131	0.86375957		
+	0.1132	0.85191465		
+	0.1133	0.84765797		
+	0.1134	0.84858168		
+	0.1135	0.85293103		
+	0.1136	0.84495729		
+	0.1137	0.86180626		
+	0.1138	0.86157634		
+	0.1139	0.85724069		
+	0.114	0.87948921		
+	0.1141	0.89038712		
+	0.1142	0.90338852		
+	0.1143	0.90908383		
+	0.1144	0.9220215		
+	0.1145	0.92860207		
+	0.1146	0.92313371		
+	0.1147	0.92724267		
+	0.1148	0.92756106		
+	0.1149	0.93823677		
+	0.115	0.95001542		
+	0.1151	0.94129994		
+	0.1152	0.94274019		
+	0.1153	0.94825007		
+	0.1154	0.95764009		
+	0.1155	0.95248295		
+	0.1156	0.96620701		
+	0.1157	0.96096638		
+	0.1158	0.96086362		
+	0.1159	0.96499763		
+	0.116	0.9545609		
+	0.1161	0.96056063		
+	0.1162	0.96122151		
+	0.1163	0.9485824		
+	0.1164	0.94730362		
+	0.1165	0.94520172		
+	0.1166	0.95446442		
+	0.1167	0.9575194		
+	0.1168	0.97364595		
+	0.1169	0.96514939		
+	0.117	0.9851014		
+	0.1171	1.0034057		
+	0.1172	1.0040582		
+	0.1173	1.0138284		
+	0.1174	1.0001355		
+	0.1175	1.0128783		
+	0.1176	1.0006127		
+	0.1177	1.0164459		
+	0.1178	1.0122218		
+	0.1179	0.99457262		
+	0.118	1.0062748		
+	0.1181	1.0019937		
+	0.1182	1.0028522		
+	0.1183	0.99907868		
+	0.1184	0.98190701		
+	0.1185	0.98269884		
+	0.1186	0.97130706		
+	0.1187	0.97105558		
+	0.1188	0.97393351		
+	0.1189	0.96035035		
+	0.119	0.95661878		
+	0.1191	0.9596243		
+	0.1192	0.95647481		
+	0.1193	0.96855807		
+	0.1194	0.96454646		
+	0.1195	0.95773058		
+	0.1196	0.97188228		
+	0.1197	0.96822353		
+	0.1198	0.97866808		
+	0.1199	0.98841043		
+	0.12	0.99564774		
+	0.1201	1.0002274		
+	0.1202	1.0047563		
+	0.1203	1.0175155		
+	0.1204	1.0154286		
+	0.1205	1.0163638		
+	0.1206	0.99609959		
+	0.1207	0.99588576		
+	0.1208	1.0031606		
+	0.1209	0.99155578		
+	0.121	0.98559819		
+	0.1211	0.96537118		
+	0.1212	0.94746663		
+	0.1213	0.93319676		
+	0.1214	0.92551242		
+	0.1215	0.91760129		
+	0.1216	0.91537875		
+	0.1217	0.91214876		
+	0.1218	0.88812713		
+	0.1219	0.89217698		
+	0.122	0.89101245		
+	0.1221	0.86764241		
+	0.1222	0.86825296		
+	0.1223	0.87670142		
+	0.1224	0.8655865		
+	0.1225	0.86496635		
+	0.1226	0.85680222		
+	0.1227	0.87023771		
+	0.1228	0.8785361		
+	0.1229	0.88538331		
+	0.123	0.90019366		
+	0.1231	0.90459968		
+	0.1232	0.89293169		
+	0.1233	0.89427402		
+	0.1234	0.89586277		
+	0.1235	0.89467111		
+	0.1236	0.90015336		
+	0.1237	0.89582765		
+	0.1238	0.88705508		
+	0.1239	0.89226638		
+	0.124	0.88706145		
+	0.1241	0.87751602		
+	0.1242	0.87055363		
+	0.1243	0.863671		
+	0.1244	0.85560065		
+	0.1245	0.85389751		
+	0.1246	0.85576792		
+	0.1247	0.84783063		
+	0.1248	0.8496618		
+	0.1249	0.84634642		
+	0.125	0.83792999		
+	0.1251	0.84062051		
+	0.1252	0.84333725		
+	0.1253	0.84559549		
+	0.1254	0.85288841		
+	0.1255	0.84729374		
+	0.1256	0.86179295		
+	0.1257	0.87042116		
+	0.1258	0.8780241		
+	0.1259	0.88331117		
+	0.126	0.89442418		
+	0.1261	0.89908169		
+	0.1262	0.88578802		
+	0.1263	0.89585585		
+	0.1264	0.89081411		
+	0.1265	0.89244751		
+	0.1266	0.88539491		
+	0.1267	0.89221461		
+	0.1268	0.87589658		
+	0.1269	0.87137483		
+	0.127	0.880487		
+	0.1271	0.8805949		
+	0.1272	0.86909579		
+	0.1273	0.86990846		
+	0.1274	0.86010299		
+	0.1275	0.86078241		
+	0.1276	0.85676397		
+	0.1277	0.85901065		
+	0.1278	0.85243071		
+	0.1279	0.8451604		
+	0.128	0.84458187		
+	0.1281	0.8464142		
+	0.1282	0.84863307		
+	0.1283	0.83494537		
+	0.1284	0.85415156		
+	0.1285	0.85876357		
+	0.1286	0.87029622		
+	0.1287	0.87697967		
+	0.1288	0.88468121		
+	0.1289	0.88715643		
+	0.129	0.89690602		
+	0.1291	0.89204119		
+	0.1292	0.88906636		
+	0.1293	0.89670531		
+	0.1294	0.89973744		
+	0.1295	0.88022556		
+	0.1296	0.88669152		
+	0.1297	0.87957077		
+	0.1298	0.88427289		
+	0.1299	0.88449605		
+	0.13	0.8717567		
+	0.1301	0.87311934		
+	0.1302	0.87382481		
+	0.1303	0.876095		
+	0.1304	0.86905336		
+	0.1305	0.85668198		
+	0.1306	0.85783984		
+	0.1307	0.87670514		
+	0.1308	0.87038803		
+	0.1309	0.87699232		
+	0.131	0.88527388		
+	0.1311	0.87586139		
+	0.1312	0.89474708		
+	0.1313	0.89532468		
+	0.1314	0.91546659		
+	0.1315	0.9300665		
+	0.1316	0.94042402		
+	0.1317	0.9465874		
+	0.1318	0.96812125		
+	0.1319	0.97636766		
+	0.132	0.97600905		
+	0.1321	0.98069804		
+	0.1322	0.99499507		
+	0.1323	0.9895055		
+	0.1324	0.99399579		
+	0.1325	0.99643631		
+	0.1326	0.98168543		
+	0.1327	0.97390884		
+	0.1328	0.97353967		
+	0.1329	0.97116095		
+	0.133	0.9735709		
+	0.1331	0.96127325		
+	0.1332	0.97417221		
+	0.1333	0.9565358		
+	0.1334	0.95581625		
+	0.1335	0.95182745		
+	0.1336	0.95432944		
+	0.1337	0.96506427		
+	0.1338	0.96013325		
+	0.1339	0.95301699		
+	0.134	0.95022177		
+	0.1341	0.95541635		
+	0.1342	0.95286374		
+	0.1343	0.95983477		
+	0.1344	0.96147723		
+	0.1345	0.98101913		
+	0.1346	0.98836388		
+	0.1347	0.99795654		
+	0.1348	1.0051541		
+	0.1349	1.0049452		
+	0.135	1.0107872		
+	0.1351	1.0111318		
+	0.1352	1.0053808		
+	0.1353	0.99415158		
+	0.1354	0.99669913		
+	0.1355	0.99329193		
+	0.1356	0.99634883		
+	0.1357	0.99726801		
+	0.1358	0.98176881		
+	0.1359	0.97839263		
+	0.136	0.97487203		
+	0.1361	0.98201289		
+	0.1362	0.96583439		
+	0.1363	0.96349516		
+	0.1364	0.95400857		
+	0.1365	0.95450542		
+	0.1366	0.94912207		
+	0.1367	0.95102826		
+	0.1368	0.94347424		
+	0.1369	0.95131333		
+	0.137	0.95245614		
+	0.1371	0.94637217		
+	0.1372	0.94565887		
+	0.1373	0.94252912		
+	0.1374	0.94598274		
+	0.1375	0.9437063		
+	0.1376	0.95749096		
+	0.1377	0.95246632		
+	0.1378	0.94624866		
+	0.1379	0.9419611		
+	0.138	0.9303728		
+	0.1381	0.92176298		
+	0.1382	0.91754366		
+	0.1383	0.91436207		
+	0.1384	0.90876059		
+	0.1385	0.90028161		
+	0.1386	0.8956743		
+	0.1387	0.88569886		
+	0.1388	0.88386625		
+	0.1389	0.88132749		
+	0.139	0.8616126		
+	0.1391	0.85531741		
+	0.1392	0.85427479		
+	0.1393	0.84931481		
+	0.1394	0.84709565		
+	0.1395	0.83583776		
+	0.1396	0.84133264		
+	0.1397	0.83096655		
+	0.1398	0.84115102		
+	0.1399	0.84167578		
+	0.14	0.83518103		
+	0.1401	0.83459339		
+	0.1402	0.85203831		
+	0.1403	0.85349988		
+	0.1404	0.86256349		
+	0.1405	0.87305385		
+	0.1406	0.8779057		
+	0.1407	0.87870758		
+	0.1408	0.8857894		
+	0.1409	0.88575693		
+	0.141	0.87599161		
+	0.1411	0.88702375		
+	0.1412	0.87116916		
+	0.1413	0.88292551		
+	0.1414	0.8674676		
+	0.1415	0.87849762		
+	0.1416	0.87421409		
+	0.1417	0.85673578		
+	0.1418	0.86031562		
+	0.1419	0.85652843		
+	0.142	0.8616933		
+	0.1421	0.84197576		
+	0.1422	0.83577451		
+	0.1423	0.83355781		
+	0.1424	0.84164636		
+	0.1425	0.83159163		
+	0.1426	0.83028438		
+	0.1427	0.82658414		
+	0.1428	0.8258147		
+	0.1429	0.83488119		
+	0.143	0.8390222		
+	0.1431	0.83889795		
+	0.1432	0.84705388		
+	0.1433	0.86363643		
+	0.1434	0.8629931		
+	0.1435	0.8860291		
+	0.1436	0.88734728		
+	0.1437	0.87801076		
+	0.1438	0.88389513		
+	0.1439	0.88023521		
+	0.144	0.8722192		
+	0.1441	0.87970972		
+	0.1442	0.8868228		
+	0.1443	0.87654351		
+	0.1444	0.8626208		
+	0.1445	0.87070062		
+	0.1446	0.86766191		
+	0.1447	0.85994919		
+	0.1448	0.8587102		
+	0.1449	0.85631336		
+	0.145	0.85229106		
+	0.1451	0.84702355		
+	0.1452	0.83377481		
+	0.1453	0.84897551		
+	0.1454	0.82925517		
+	0.1455	0.8434522		
+	0.1456	0.84447069		
+	0.1457	0.82374609		
+	0.1458	0.83677438		
+	0.1459	0.83383523		
+	0.146	0.84363489		
+	0.1461	0.84447272		
+	0.1462	0.85831115		
+	0.1463	0.88023064		
+	0.1464	0.87639471		
+	0.1465	0.88222553		
+	0.1466	0.90142626		
+	0.1467	0.8989444		
+	0.1468	0.9024676		
+	0.1469	0.9069272		
+	0.147	0.89371739		
+	0.1471	0.89311636		
+	0.1472	0.89663268		
+	0.1473	0.90931054		
+	0.1474	0.91168676		
+	0.1475	0.91424315		
+	0.1476	0.90449141		
+	0.1477	0.92390249		
+	0.1478	0.91296375		
+	0.1479	0.91192691		
+	0.148	0.92395398		
+	0.1481	0.91539115		
+	0.1482	0.93121295		
+	0.1483	0.92014374		
+	0.1484	0.92260129		
+	0.1485	0.92797376		
+	0.1486	0.93933169		
+	0.1487	0.94062332		
+	0.1488	0.92447372		
+	0.1489	0.93796674		
+	0.149	0.93811233		
+	0.1491	0.96687838		
+	0.1492	0.96932449		
+	0.1493	0.97273491		
+	0.1494	0.99380512		
+	0.1495	0.98223561		
+	0.1496	0.98845226		
+	0.1497	0.98405146		
+	0.1498	0.99608527		
+	0.1499	0.99498531		
+	0.15	0.97768401		
+	0.1501	0.98461206		
+	0.1502	0.97549537		
+	0.1503	0.97459173		
+	0.1504	0.97725608		
+	0.1505	0.96409021		
+	0.1506	0.97315743		
+	0.1507	0.96655008		
+	0.1508	0.95234336		
+	0.1509	0.96505751		
+	0.151	0.94621904		
+	0.1511	0.94931648		
+	0.1512	0.95263134		
+	0.1513	0.95435323		
+	0.1514	0.93552449		
+	0.1515	0.93298821		
+	0.1516	0.93604422		
+	0.1517	0.93961022		
+	0.1518	0.94355018		
+	0.1519	0.96121655		
+	0.152	0.96712655		
+	0.1521	0.96580506		
+	0.1522	0.97399686		
+	0.1523	0.98944508		
+	0.1524	0.99913506		
+	0.1525	0.99057135		
+	0.1526	0.98972403		
+	0.1527	0.98343196		
+	0.1528	0.98022578		
+	0.1529	0.99223309		
+	0.153	0.98948298		
+	0.1531	0.9841798		
+	0.1532	0.98147796		
+	0.1533	0.97850681		
+	0.1534	0.961368		
+	0.1535	0.94868798		
+	0.1536	0.94544739		
+	0.1537	0.93288568		
+	0.1538	0.90813269		
+	0.1539	0.90075838		
+	0.154	0.90044248		
+	0.1541	0.88406374		
+	0.1542	0.88241033		
+	0.1543	0.87797073		
+	0.1544	0.87014072		
+	0.1545	0.85398686		
+	0.1546	0.86816462		
+	0.1547	0.85109855		
+	0.1548	0.86719436		
+	0.1549	0.87152126		
+	0.155	0.87331009		
+	0.1551	0.87363259		
+	0.1552	0.89485842		
+	0.1553	0.89356673		
+	0.1554	0.87641859		
+	0.1555	0.88551022		
+	0.1556	0.88108036		
+	0.1557	0.8737304		
+	0.1558	0.86395145		
+	0.1559	0.86692005		
+	0.156	0.86584385		
+	0.1561	0.86951146		
+	0.1562	0.86686607		
+	0.1563	0.86377998		
+	0.1564	0.84297441		
+	0.1565	0.84361465		
+	0.1566	0.85001456		
+	0.1567	0.82956854		
+	0.1568	0.83455092		
+	0.1569	0.83705759		
+	0.157	0.82982262		
+	0.1571	0.82703383		
+	0.1572	0.82337832		
+	0.1573	0.83309544		
+	0.1574	0.81590923		
+	0.1575	0.81718451		
+	0.1576	0.82932272		
+	0.1577	0.82831287		
+	0.1578	0.8470732		
+	0.1579	0.84032722		
+	0.158	0.85982433		
+	0.1581	0.86282896		
+	0.1582	0.8752929		
+	0.1583	0.87260648		
+	0.1584	0.86877295		
+	0.1585	0.87398234		
+	0.1586	0.86907814		
+	0.1587	0.85972796		
+	0.1588	0.8617113		
+	0.1589	0.85823101		
+	0.159	0.86589656		
+	0.1591	0.85617656		
+	0.1592	0.86336009		
+	0.1593	0.8541		
+	0.1594	0.84522593		
+	0.1595	0.84633811		
+	0.1596	0.84323779		
+	0.1597	0.82817621		
+	0.1598	0.82650515		
+	0.1599	0.83791111		
+	0.16	0.82848127		
+	0.1601	0.81688744		
+	0.1602	0.82793201		
+	0.1603	0.82809056		
+	0.1604	0.81669529		
+	0.1605	0.81389604		
+	0.1606	0.82501088		
+	0.1607	0.82935885		
+	0.1608	0.83870222		
+	0.1609	0.86092552		
+	0.161	0.85970756		
+	0.1611	0.86171742		
+	0.1612	0.87605922		
+	0.1613	0.8737332		
+	0.1614	0.86629583		
+	0.1615	0.86814254		
+	0.1616	0.86924918		
+	0.1617	0.87080524		
+	0.1618	0.85856779		
+	0.1619	0.87165948		
+	0.162	0.85095327		
+	0.1621	0.85729281		
+	0.1622	0.84213548		
+	0.1623	0.85660415		
+	0.1624	0.84067315		
+	0.1625	0.84097793		
+	0.1626	0.84672762		
+	0.1627	0.83511054		
+	0.1628	0.83767307		
+	0.1629	0.83051983		
+	0.163	0.83651152		
+	0.1631	0.84324401		
+	0.1632	0.84871334		
+	0.1633	0.84980971		
+	0.1634	0.84986392		
+	0.1635	0.85615243		
+	0.1636	0.86681964		
+	0.1637	0.87695345		
+	0.1638	0.90468929		
+	0.1639	0.92133547		
+	0.164	0.92196747		
+	0.1641	0.93364746		
+	0.1642	0.94650959		
+	0.1643	0.95336073		
+	0.1644	0.94767525		
+	0.1645	0.95105874		
+	0.1646	0.9498333		
+	0.1647	0.96597942		
+	0.1648	0.95142989		
+	0.1649	0.95500443		
+	0.165	0.94716273		
+	0.1651	0.9534483		
+	0.1652	0.9554155		
+	0.1653	0.95413014		
+	0.1654	0.94492501		
+	0.1655	0.93155138		
+	0.1656	0.93956981		
+	0.1657	0.93859519		
+	0.1658	0.92921398		
+	0.1659	0.92254327		
+	0.166	0.93632551		
+	0.1661	0.9291106		
+	0.1662	0.92607262		
+	0.1663	0.9224375		
+	0.1664	0.93864609		
+	0.1665	0.94360548		
+	0.1666	0.94650386		
+	0.1667	0.96150594		
+	0.1668	0.96975764		
+	0.1669	0.97829855		
+	0.167	0.9824415		
+	0.1671	0.98941923		
+	0.1672	0.98566153		
+	0.1673	0.97749585		
+	0.1674	0.98183805		
+	0.1675	0.9681756		
+	0.1676	0.97392807		
+	0.1677	0.98243118		
+	0.1678	0.97333838		
+	0.1679	0.97320658		
+	0.168	0.96783436		
+	0.1681	0.95551205		
+	0.1682	0.95219674		
+	0.1683	0.94174868		
+	0.1684	0.94513895		
+	0.1685	0.94537306		
+	0.1686	0.93116073		
+	0.1687	0.9360817		
+	0.1688	0.92807132		
+	0.1689	0.92805568		
+	0.169	0.92432543		
+	0.1691	0.93278171		
+	0.1692	0.93883176		
+	0.1693	0.93225917		
+	0.1694	0.93137029		
+	0.1695	0.93307991		
+	0.1696	0.9594042		
+	0.1697	0.94923701		
+	0.1698	0.96809974		
+	0.1699	0.950353		
+	0.17	0.95297763		
+	0.1701	0.94359494		
+	0.1702	0.93649749		
+	0.1703	0.92205309		
+	0.1704	0.91883452		
+	0.1705	0.90841179		
+	0.1706	0.90951334		
+	0.1707	0.88858774		
+	0.1708	0.88698309		
+	0.1709	0.87018051		
+	0.171	0.8764923		
+	0.1711	0.86674792		
+	0.1712	0.86151369		
+	0.1713	0.84711463		
+	0.1714	0.83485709		
+	0.1715	0.84424896		
+	0.1716	0.82890557		
+	0.1717	0.82620086		
+	0.1718	0.83167602		
+	0.1719	0.8128626		
+	0.172	0.81826091		
+	0.1721	0.82103425		
+	0.1722	0.81365033		
+	0.1723	0.81873659		
+	0.1724	0.82085382		
+	0.1725	0.83374626		
+	0.1726	0.85238879		
+	0.1727	0.85312977		
+	0.1728	0.86487366		
+	0.1729	0.85841276		
+	0.173	0.87032129		
+	0.1731	0.8623362		
+	0.1732	0.86547496		
+	0.1733	0.85404911		
+	0.1734	0.85429785		
+	0.1735	0.86299895		
+	0.1736	0.84397335		
+	0.1737	0.84384245		
+	0.1738	0.84599858		
+	0.1739	0.84573507		
+	0.174	0.84584348		
+	0.1741	0.84142141		
+	0.1742	0.83828939		
+	0.1743	0.82157941		
+	0.1744	0.83119226		
+	0.1745	0.80991444		
+	0.1746	0.8167318		
+	0.1747	0.81636856		
+	0.1748	0.81667466		
+	0.1749	0.81719736		
+	0.175	0.81014505		
+	0.1751	0.80215641		
+	0.1752	0.81586232		
+	0.1753	0.8308756		
+	0.1754	0.8405025		
+	0.1755	0.84393005		
+	0.1756	0.85822261		
+	0.1757	0.86943062		
+	0.1758	0.85367373		
+	0.1759	0.86647853		
+	0.176	0.87166613		
+	0.1761	0.85653946		
+	0.1762	0.85990391		
+	0.1763	0.85417557		
+	0.1764	0.84610378		
+	0.1765	0.84847513		
+	0.1766	0.84256036		
+	0.1767	0.83771313		
+	0.1768	0.83175422		
+	0.1769	0.83555389		
+	0.177	0.8355314		
+	0.1771	0.83584187		
+	0.1772	0.82169274		
+	0.1773	0.82252577		
+	0.1774	0.82160058		
+	0.1775	0.82534171		
+	0.1776	0.82146603		
+	0.1777	0.81452446		
+	0.1778	0.8032786		
+	0.1779	0.81777747		
+	0.178	0.81611348		
+	0.1781	0.81268424		
+	0.1782	0.828693		
+	0.1783	0.82699591		
+	0.1784	0.84196782		
+	0.1785	0.85660564		
+	0.1786	0.85918885		
+	0.1787	0.86791		
+	0.1788	0.86763788		
+	0.1789	0.86581815		
+	0.179	0.85599954		
+	0.1791	0.86696334		
+	0.1792	0.85746792		
+	0.1793	0.86061283		
+	0.1794	0.87398512		
+	0.1795	0.87046775		
+	0.1796	0.86497236		
+	0.1797	0.87455088		
+	0.1798	0.86313375		
+	0.1799	0.87345287		
+	0.18	0.8766108		
+	0.1801	0.8735995		
+	0.1802	0.87480398		
+	0.1803	0.88736746		
+	0.1804	0.87664619		
+	0.1805	0.89171837		
+	0.1806	0.89413719		
+	0.1807	0.89502673		
+	0.1808	0.90752202		
+	0.1809	0.91213241		
+	0.181	0.90276135		
+	0.1811	0.91049548		
+	0.1812	0.92022708		
+	0.1813	0.93050045		
+	0.1814	0.9555712		
+	0.1815	0.95995495		
+	0.1816	0.96106057		
+	0.1817	0.96904925		
+	0.1818	0.9672497		
+	0.1819	0.96968482		
+	0.182	0.96075194		
+	0.1821	0.96749485		
+	0.1822	0.95943118		
+	0.1823	0.95682923		
+	0.1824	0.94954244		
+	0.1825	0.94587833		
+	0.1826	0.95043062		
+	0.1827	0.93738602		
+	0.1828	0.949155		
+	0.1829	0.94068021		
+	0.183	0.93244175		
+	0.1831	0.93512691		
+	0.1832	0.93762102		
+	0.1833	0.92166614		
+	0.1834	0.91730385		
+	0.1835	0.91776674		
+	0.1836	0.92901555		
+	0.1837	0.91991586		
+	0.1838	0.91524822		
+	0.1839	0.91312939		
+	0.184	0.92081102		
+	0.1841	0.93982925		
+	0.1842	0.93977143		
+	0.1843	0.95736933		
+	0.1844	0.96374511		
+	0.1845	0.9718438		
+	0.1846	0.97371836		
+	0.1847	0.97193359		
+	0.1848	0.96194717		
+	0.1849	0.97224343		
+	0.185	0.96201446		
+	0.1851	0.96238156		
+	0.1852	0.96139331		
+	0.1853	0.95080328		
+	0.1854	0.95344523		
+	0.1855	0.95934101		
+	0.1856	0.95496132		
+	0.1857	0.93243181		
+	0.1858	0.92970749		
+	0.1859	0.93146612		
+	0.186	0.92611678		
+	0.1861	0.91114104		
+	0.1862	0.90241943		
+	0.1863	0.88511656		
+	0.1864	0.87610057		
+	0.1865	0.88316118		
+	0.1866	0.86607822		
+	0.1867	0.84992382		
+	0.1868	0.86230265		
+	0.1869	0.84669856		
+	0.187	0.85679534		
+	0.1871	0.86034086		
+	0.1872	0.87439128		
+	0.1873	0.88461841		
+	0.1874	0.88290011		
+	0.1875	0.88104939		
+	0.1876	0.87481858		
+	0.1877	0.87641587		
+	0.1878	0.8635625		
+	0.1879	0.86968427		
+	0.188	0.85175741		
+	0.1881	0.85800753		
+	0.1882	0.85747405		
+	0.1883	0.83774714		
+	0.1884	0.82927598		
+	0.1885	0.84122738		
+	0.1886	0.82278082		
+	0.1887	0.82423129		
+	0.1888	0.8237352		
+	0.1889	0.81960705		
+	0.189	0.81277737		
+	0.1891	0.81431151		
+	0.1892	0.81074469		
+	0.1893	0.80064553		
+	0.1894	0.81293834		
+	0.1895	0.80059357		
+	0.1896	0.80226382		
+	0.1897	0.79729924		
+	0.1898	0.80737621		
+	0.1899	0.81325913		
+	0.19	0.81516499		
+	0.1901	0.83419682		
+	0.1902	0.8487807		
+	0.1903	0.84510508		
+	0.1904	0.84259803		
+	0.1905	0.8468928		
+	0.1906	0.84495733		
+	0.1907	0.84952666		
+	0.1908	0.84008683		
+	0.1909	0.85663958		
+	0.191	0.84888472		
+	0.1911	0.8476218		
+	0.1912	0.8321953		
+	0.1913	0.83621457		
+	0.1914	0.82698374		
+	0.1915	0.8345029		
+	0.1916	0.82322058		
+	0.1917	0.81163753		
+	0.1918	0.81993509		
+	0.1919	0.81164855		
+	0.192	0.80120477		
+	0.1921	0.80860874		
+	0.1922	0.80599034		
+	0.1923	0.80345093		
+	0.1924	0.80780258		
+	0.1925	0.80200771		
+	0.1926	0.80385784		
+	0.1927	0.81061245		
+	0.1928	0.81034525		
+	0.1929	0.81973161		
+	0.193	0.83674911		
+	0.1931	0.84125375		
+	0.1932	0.8538518		
+	0.1933	0.84862363		
+	0.1934	0.86133765		
+	0.1935	0.84719787		
+	0.1936	0.85333903		
+	0.1937	0.85096878		
+	0.1938	0.84704865		
+	0.1939	0.83615419		
+	0.194	0.84478381		
+	0.1941	0.83202012		
+	0.1942	0.82810944		
+	0.1943	0.84023392		
+	0.1944	0.82746454		
+	0.1945	0.82785464		
+	0.1946	0.82053933		
+	0.1947	0.81978458		
+	0.1948	0.80445564		
+	0.1949	0.80742583		
+	0.195	0.81231062		
+	0.1951	0.80835529		
+	0.1952	0.80549341		
+	0.1953	0.80484216		
+	0.1954	0.80234472		
+	0.1955	0.80910667		
+	0.1956	0.81811547		
+	0.1957	0.82642847		
+	0.1958	0.83442369		
+	0.1959	0.85577365		
+	0.196	0.85930708		
+	0.1961	0.87446631		
+	0.1962	0.89107658		
+	0.1963	0.89390853		
+	0.1964	0.90741947		
+	0.1965	0.90936999		
+	0.1966	0.90969646		
+	0.1967	0.90484829		
+	0.1968	0.9270459		
+	0.1969	0.91504508		
+	0.197	0.92599854		
+	0.1971	0.92400991		
+	0.1972	0.92919984		
+	0.1973	0.91888106		
+	0.1974	0.92800021		
+	0.1975	0.91277128		
+	0.1976	0.92521596		
+	0.1977	0.90513612		
+	0.1978	0.91546742		
+	0.1979	0.91167234		
+	0.198	0.90098422		
+	0.1981	0.91416123		
+	0.1982	0.9079211		
+	0.1983	0.89528712		
+	0.1984	0.91359625		
+	0.1985	0.91362876		
+	0.1986	0.91080795		
+	0.1987	0.91701139		
+	0.1988	0.93310671		
+	0.1989	0.94542105		
+	0.199	0.94959662		
+	0.1991	0.95198393		
+	0.1992	0.9587513		
+	0.1993	0.96706499		
+	0.1994	0.95666641		
+	0.1995	0.95866186		
+	0.1996	0.95550924		
+	0.1997	0.94719292		
+	0.1998	0.95861105		
+	0.1999	0.94748332		
+	0.2	0.94361814		
+	0.2001	0.94140392		
+	0.2002	0.93783727		
+	0.2003	0.93275506		
+	0.2004	0.92661982		
+	0.2005	0.93612927		
+	0.2006	0.92864443		
+	0.2007	0.92884099		
+	0.2008	0.90894544		
+	0.2009	0.91811164		
+	0.201	0.9086156		
+	0.2011	0.91418995		
+	0.2012	0.91748088		
+	0.2013	0.91579192		
+	0.2014	0.91638691		
+	0.2015	0.90570407		
+	0.2016	0.92508202		
+	0.2017	0.93281028		
+	0.2018	0.9344626		
+	0.2019	0.95800019		
+	0.202	0.95063627		
+	0.2021	0.94690637		
+	0.2022	0.94675733		
+	0.2023	0.94690135		
+	0.2024	0.93630447		
+	0.2025	0.93227808		
+	0.2026	0.92527762		
+	0.2027	0.9088977		
+	0.2028	0.90532414		
+	0.2029	0.89962776		
+	0.203	0.88745603		
+	0.2031	0.87526522		
+	0.2032	0.86847735		
+	0.2033	0.8509887		
+	0.2034	0.84716192		
+	0.2035	0.83656263		
+	0.2036	0.83739658		
+	0.2037	0.82949569		
+	0.2038	0.81611549		
+	0.2039	0.80842741		
+	0.204	0.81028945		
+	0.2041	0.79985913		
+	0.2042	0.80676428		
+	0.2043	0.79323091		
+	0.2044	0.7984423		
+	0.2045	0.81045263		
+	0.2046	0.8054725		
+	0.2047	0.8221023		
+	0.2048	0.8411093		
+	0.2049	0.84519345		
+	0.205	0.83587248		
+	0.2051	0.84913576		
+	0.2052	0.85064115		
+	0.2053	0.83262534		
+	0.2054	0.84500075		
+	0.2055	0.84657872		
+	0.2056	0.84018655		
+	0.2057	0.83664347		
+	0.2058	0.82114655		
+	0.2059	0.8189266		
+	0.206	0.82684122		
+	0.2061	0.82589242		
+	0.2062	0.81340164		
+	0.2063	0.81806154		
+	0.2064	0.8105014		
+	0.2065	0.79568251		
+	0.2066	0.80433549		
+	0.2067	0.79758658		
+	0.2068	0.80047319		
+	0.2069	0.79865565		
+	0.207	0.79111144		
+	0.2071	0.78455527		
+	0.2072	0.79434657		
+	0.2073	0.79826514		
+	0.2074	0.78920063		
+	0.2075	0.80975906		
+	0.2076	0.8246757		
+	0.2077	0.82140206		
+	0.2078	0.83979006		
+	0.2079	0.84337501		
+	0.208	0.85285004		
+	0.2081	0.84278772		
+	0.2082	0.84275223		
+	0.2083	0.83343867		
+	0.2084	0.83278237		
+	0.2085	0.83146875		
+	0.2086	0.84121243		
+	0.2087	0.82421192		
+	0.2088	0.82145774		
+	0.2089	0.82964108		
+	0.209	0.8146301		
+	0.2091	0.81430775		
+	0.2092	0.8083464		
+	0.2093	0.80113033		
+	0.2094	0.81113381		
+	0.2095	0.79460476		
+	0.2096	0.80381247		
+	0.2097	0.80598808		
+	0.2098	0.79829863		
+	0.2099	0.7975013		
+	0.21	0.79341482		
+	0.2101	0.78711369		
+	0.2102	0.78485551		
+	0.2103	0.79784663		
+	0.2104	0.80166718		
+	0.2105	0.82313277		
+	0.2106	0.82437127		
+	0.2107	0.84211186		
+	0.2108	0.84742928		
+	0.2109	0.83641123		
+	0.211	0.8464829		
+	0.2111	0.84704173		
+	0.2112	0.8443986		
+	0.2113	0.84412413		
+	0.2114	0.83799125		
+	0.2115	0.82764058		
+	0.2116	0.82640659		
+	0.2117	0.83545053		
+	0.2118	0.83376986		
+	0.2119	0.8238891		
+	0.212	0.83084824		
+	0.2121	0.8351752		
+	0.2122	0.82941218		
+	0.2123	0.84073608		
+	0.2124	0.8412473		
+	0.2125	0.84594491		
+	0.2126	0.83141753		
+	0.2127	0.8495859		
+	0.2128	0.84979833		
+	0.2129	0.84834267		
+	0.213	0.86676859		
+	0.2131	0.86334241		
+	0.2132	0.87333415		
+	0.2133	0.89006689		
+	0.2134	0.9059871		
+	0.2135	0.90939002		
+	0.2136	0.93613312		
+	0.2137	0.927387		
+	0.2138	0.94561376		
+	0.2139	0.95292756		
+	0.214	0.95313541		
+	0.2141	0.93921183		
+	0.2142	0.935933		
+	0.2143	0.93305357		
+	0.2144	0.94394754		
+	0.2145	0.92677042		
+	0.2146	0.92944776		
+	0.2147	0.92087541		
+	0.2148	0.93389393		
+	0.2149	0.92604683		
+	0.215	0.92369891		
+	0.2151	0.91432192		
+	0.2152	0.91447501		
+	0.2153	0.91127043		
+	0.2154	0.89988261		
+	0.2155	0.91040944		
+	0.2156	0.90623677		
+	0.2157	0.90717343		
+	0.2158	0.9015931		
+	0.2159	0.90365972		
+	0.216	0.90757234		
+	0.2161	0.90966535		
+	0.2162	0.91057429		
+	0.2163	0.92490755		
+	0.2164	0.9369037		
+	0.2165	0.93977704		
+	0.2166	0.94409296		
+	0.2167	0.95831545		
+	0.2168	0.96198526		
+	0.2169	0.96251706		
+	0.217	0.95094617		
+	0.2171	0.95067285		
+	0.2172	0.95499137		
+	0.2173	0.95440425		
+	0.2174	0.95218679		
+	0.2175	0.9450745		
+	0.2176	0.94263846		
+	0.2177	0.93600287		
+	0.2178	0.93851541		
+	0.2179	0.9339802		
+	0.218	0.92379877		
+	0.2181	0.92363817		
+	0.2182	0.91274448		
+	0.2183	0.91227032		
+	0.2184	0.90493795		
+	0.2185	0.9054429		
+	0.2186	0.88823013		
+	0.2187	0.88225867		
+	0.2188	0.87018165		
+	0.2189	0.86264038		
+	0.219	0.86382022		
+	0.2191	0.85740544		
+	0.2192	0.85575367		
+	0.2193	0.87634585		
+	0.2194	0.8838637		
+	0.2195	0.88585528		
+	0.2196	0.88662672		
+	0.2197	0.87329874		
+	0.2198	0.87118302		
+	0.2199	0.85967599		
+	0.22	0.86606687		
+	0.2201	0.85683414		
+	0.2202	0.84591905		
+	0.2203	0.85175389		
+	0.2204	0.84821226		
+	0.2205	0.83689393		
+	0.2206	0.82174021		
+	0.2207	0.81678677		
+	0.2208	0.81467305		
+	0.2209	0.8029601		
+	0.221	0.79572282		
+	0.2211	0.79749943		
+	0.2212	0.7866808		
+	0.2213	0.80133967		
+	0.2214	0.79813405		
+	0.2215	0.79708874		
+	0.2216	0.7872825		
+	0.2217	0.79456286		
+	0.2218	0.78259066		
+	0.2219	0.77821517		
+	0.222	0.7930902		
+	0.2221	0.79942595		
+	0.2222	0.8163156		
+	0.2223	0.82488215		
+	0.2224	0.82433718		
+	0.2225	0.82680515		
+	0.2226	0.83972513		
+	0.2227	0.83350395		
+	0.2228	0.83708704		
+	0.2229	0.83043297		
+	0.223	0.82734795		
+	0.2231	0.83095999		
+	0.2232	0.82144486		
+	0.2233	0.81804562		
+	0.2234	0.82616546		
+	0.2235	0.82008718		
+	0.2236	0.82013339		
+	0.2237	0.80066337		
+	0.2238	0.80732727		
+	0.2239	0.79906703		
+	0.224	0.7935783		
+	0.2241	0.7874804		
+	0.2242	0.7933762		
+	0.2243	0.78908378		
+	0.2244	0.78901255		
+	0.2245	0.79470387		
+	0.2246	0.77832823		
+	0.2247	0.78621801		
+	0.2248	0.77775805		
+	0.2249	0.79314067		
+	0.225	0.79859547		
+	0.2251	0.80812441		
+	0.2252	0.82464336		
+	0.2253	0.82578148		
+	0.2254	0.82526138		
+	0.2255	0.83581399		
+	0.2256	0.83397579		
+	0.2257	0.8287265		
+	0.2258	0.83681741		
+	0.2259	0.83669192		
+	0.226	0.83154968		
+	0.2261	0.82110333		
+	0.2262	0.83419786		
+	0.2263	0.81360933		
+	0.2264	0.81436436		
+	0.2265	0.8089145		
+	0.2266	0.81710405		
+	0.2267	0.81127503		
+	0.2268	0.80590054		
+	0.2269	0.80958576		
+	0.227	0.80367386		
+	0.2271	0.79405286		
+	0.2272	0.79590769		
+	0.2273	0.78317198		
+	0.2274	0.79824648		
+	0.2275	0.78053388		
+	0.2276	0.78378299		
+	0.2277	0.79182563		
+	0.2278	0.78511504		
+	0.2279	0.79083667		
+	0.228	0.81567632		
+	0.2281	0.81629183		
+	0.2282	0.82626983		
+	0.2283	0.84223462		
+	0.2284	0.86201686		
+	0.2285	0.85879079		
+	0.2286	0.86734248		
+	0.2287	0.86561477		
+	0.2288	0.8805524		
+	0.2289	0.88284584		
+	0.229	0.87620387		
+	0.2291	0.87582591		
+	0.2292	0.88777297		
+	0.2293	0.88064203		
+	0.2294	0.89420354		
+	0.2295	0.89144104		
+	0.2296	0.90181346		
+	0.2297	0.90177261		
+	0.2298	0.89827316		
+	0.2299	0.8865894		
+	0.23	0.89725507		
+	0.2301	0.89062743		
+	0.2302	0.89922036		
+	0.2303	0.88588138		
+	0.2304	0.88051417		
+	0.2305	0.88300694		
+	0.2306	0.88081248		
+	0.2307	0.89320087		
+	0.2308	0.89569259		
+	0.2309	0.8982219		
+	0.231	0.92500076		
+	0.2311	0.92420629		
+	0.2312	0.93933886		
+	0.2313	0.93632603		
+	0.2314	0.9448604		
+	0.2315	0.93699236		
+	0.2316	0.93898698		
+	0.2317	0.94192186		
+	0.2318	0.93990298		
+	0.2319	0.93413271		
+	0.232	0.93548639		
+	0.2321	0.93472517		
+	0.2322	0.92666296		
+	0.2323	0.92801943		
+	0.2324	0.92386064		
+	0.2325	0.91604518		
+	0.2326	0.9185507		
+	0.2327	0.92125541		
+	0.2328	0.90703128		
+	0.2329	0.90160894		
+	0.233	0.89524963		
+	0.2331	0.91136676		
+	0.2332	0.90094769		
+	0.2333	0.8941779		
+	0.2334	0.89838927		
+	0.2335	0.88750608		
+	0.2336	0.90607342		
+	0.2337	0.90316611		
+	0.2338	0.91188157		
+	0.2339	0.92734069		
+	0.234	0.93484967		
+	0.2341	0.93441175		
+	0.2342	0.95335661		
+	0.2343	0.94766496		
+	0.2344	0.95228022		
+	0.2345	0.94422638		
+	0.2346	0.93600032		
+	0.2347	0.94366154		
+	0.2348	0.93398365		
+	0.2349	0.92933678		
+	0.235	0.92254733		
+	0.2351	0.91829418		
+	0.2352	0.89917938		
+	0.2353	0.87827222		
+	0.2354	0.88287322		
+	0.2355	0.86800753		
+	0.2356	0.84640219		
+	0.2357	0.85424638		
+	0.2358	0.84514245		
+	0.2359	0.82646844		
+	0.236	0.8325793		
+	0.2361	0.81546991		
+	0.2362	0.81805806		
+	0.2363	0.80738415		
+	0.2364	0.80637442		
+	0.2365	0.79528902		
+	0.2366	0.80129445		
+	0.2367	0.81332355		
+	0.2368	0.81978295		
+	0.2369	0.82901569		
+	0.237	0.82897768		
+	0.2371	0.84024912		
+	0.2372	0.83455297		
+	0.2373	0.83527751		
+	0.2374	0.82894159		
+	0.2375	0.82851315		
+	0.2376	0.83388993		
+	0.2377	0.82657702		
+	0.2378	0.82604898		
+	0.2379	0.82868656		
+	0.238	0.81227151		
+	0.2381	0.81846667		
+	0.2382	0.80145888		
+	0.2383	0.80081709		
+	0.2384	0.80891441		
+	0.2385	0.80462647		
+	0.2386	0.78733578		
+	0.2387	0.79298479		
+	0.2388	0.78221127		
+	0.2389	0.78426912		
+	0.239	0.78886855		
+	0.2391	0.79198454		
+	0.2392	0.77375825		
+	0.2393	0.78895176		
+	0.2394	0.77627079		
+	0.2395	0.77651524		
+	0.2396	0.79238395		
+	0.2397	0.80305813		
+	0.2398	0.80787787		
+	0.2399	0.81561745		
+	0.24	0.8264056		
+	0.2401	0.83023675		
+	0.2402	0.84180262		
+	0.2403	0.82796196		
+	0.2404	0.82246093		
+	0.2405	0.83577567		
+	0.2406	0.82743293		
+	0.2407	0.82432956		
+	0.2408	0.82478005		
+	0.2409	0.82252425		
+	0.241	0.81429902		
+	0.2411	0.81895159		
+	0.2412	0.8018362		
+	0.2413	0.79596952		
+	0.2414	0.80907044		
+	0.2415	0.79143311		
+	0.2416	0.7977615		
+	0.2417	0.79686939		
+	0.2418	0.78061368		
+	0.2419	0.79466781		
+	0.242	0.78676732		
+	0.2421	0.78494003		
+	0.2422	0.7803454		
+	0.2423	0.78485087		
+	0.2424	0.78202108		
+	0.2425	0.78940767		
+	0.2426	0.79888261		
+	0.2427	0.80314841		
+	0.2428	0.81396357		
+	0.2429	0.82535393		
+	0.243	0.83112336		
+	0.2431	0.83976709		
+	0.2432	0.8352773		
+	0.2433	0.82942722		
+	0.2434	0.82716232		
+	0.2435	0.82620971		
+	0.2436	0.83147309		
+	0.2437	0.81962587		
+	0.2438	0.8160995		
+	0.2439	0.81003587		
+	0.244	0.8128811		
+	0.2441	0.80690989		
+	0.2442	0.80170985		
+	0.2443	0.80719253		
+	0.2444	0.81081763		
+	0.2445	0.81003231		
+	0.2446	0.8002473		
+	0.2447	0.80747139		
+	0.2448	0.80248538		
+	0.2449	0.81405784		
+	0.245	0.82503928		
+	0.2451	0.81823307		
+	0.2452	0.83199702		
+	0.2453	0.82821223		
+	0.2454	0.84579761		
+	0.2455	0.85861439		
+	0.2456	0.87775132		
+	0.2457	0.89641245		
+	0.2458	0.9091001		
+	0.2459	0.92151679		
+	0.246	0.91680234		
+	0.2461	0.92024323		
+	0.2462	0.92347598		
+	0.2463	0.92559982		
+	0.2464	0.92967495		
+	0.2465	0.93449303		
+	0.2466	0.91851217		
+	0.2467	0.92634628		
+	0.2468	0.9263949		
+	0.2469	0.91315144		
+	0.247	0.91385099		
+	0.2471	0.91610276		
+	0.2472	0.91699727		
+	0.2473	0.91031497		
+	0.2474	0.90485146		
+	0.2475	0.90901216		
+	0.2476	0.90444555		
+	0.2477	0.90627823		
+	0.2478	0.89989277		
+	0.2479	0.8990016		
+	0.248	0.89826029		
+	0.2481	0.8917011		
+	0.2482	0.88935695		
+	0.2483	0.90303715		
+	0.2484	0.9037412		
+	0.2485	0.91909878		
+	0.2486	0.91777064		
+	0.2487	0.9414112		
+	0.2488	0.93411377		
+	0.2489	0.95512957		
+	0.249	0.94918847		
+	0.2491	0.94612509		
+	0.2492	0.95113121		
+	0.2493	0.94146059		
+	0.2494	0.94539988		
+	0.2495	0.9443614		
+	0.2496	0.93476918		
+	0.2497	0.93438326		
+	0.2498	0.92034351		
+	0.2499	0.91829953		
+	0.25	0.92959859		
+	0.2501	0.91628099		
+	0.2502	0.91768676		
+	0.2503	0.90692833		
+	0.2504	0.90431602		
+	0.2505	0.9121394		
+	0.2506	0.90885848		
+	0.2507	0.89180457		
+	0.2508	0.90393048		
+	0.2509	0.89659448		
+	0.251	0.88715183		
+	0.2511	0.88088499		
+	0.2512	0.89388043		
+	0.2513	0.89534697		
+	0.2514	0.89262838		
+	0.2515	0.8878036		
+	0.2516	0.8976566		
+	0.2517	0.89033199		
+	0.2518	0.89676564		
+	0.2519	0.89039453		
+	0.252	0.89083107		
+	0.2521	0.88606236		
+	0.2522	0.87278565		
+	0.2523	0.86113823		
+	0.2524	0.86278724		
+	0.2525	0.85577427		
+	0.2526	0.83915108		
+	0.2527	0.83728422		
+	0.2528	0.82897594		
+	0.2529	0.82911773		
+	0.253	0.82107049		
+	0.2531	0.81018654		
+	0.2532	0.81188629		
+	0.2533	0.79112632		
+	0.2534	0.80183009		
+	0.2535	0.782239		
+	0.2536	0.79291254		
+	0.2537	0.79111039		
+	0.2538	0.78569963		
+	0.2539	0.78716955		
+	0.254	0.77335269		
+	0.2541	0.7769684		
+	0.2542	0.79394156		
+	0.2543	0.78699371		
+	0.2544	0.8151726		
+	0.2545	0.82082422		
+	0.2546	0.82741585		
+	0.2547	0.83342219		
+	0.2548	0.82760022		
+	0.2549	0.83453863		
+	0.255	0.82291184		
+	0.2551	0.82098186		
+	0.2552	0.83127469		
+	0.2553	0.81501497		
+	0.2554	0.81900113		
+	0.2555	0.82713557		
+	0.2556	0.82307162		
+	0.2557	0.80701201		
+	0.2558	0.81129672		
+	0.2559	0.79514664		
+	0.256	0.79505692		
+	0.2561	0.79055428		
+	0.2562	0.79128213		
+	0.2563	0.78382523		
+	0.2564	0.79228684		
+	0.2565	0.77922408		
+	0.2566	0.79143334		
+	0.2567	0.77978234		
+	0.2568	0.77311744		
+	0.2569	0.78822072		
+	0.257	0.79007529		
+	0.2571	0.78259023		
+	0.2572	0.79467393		
+	0.2573	0.81162418		
+	0.2574	0.82383536		
+	0.2575	0.81887699		
+	0.2576	0.82925433		
+	0.2577	0.82913778		
+	0.2578	0.83596306		
+	0.2579	0.83257246		
+	0.258	0.82242069		
+	0.2581	0.83394352		
+	0.2582	0.82088374		
+	0.2583	0.82190495		
+	0.2584	0.81503099		
+	0.2585	0.81640843		
+	0.2586	0.80893345		
+	0.2587	0.81178429		
+	0.2588	0.79703582		
+	0.2589	0.80434146		
+	0.259	0.79925186		
+	0.2591	0.79637155		
+	0.2592	0.78667133		
+	0.2593	0.79288639		
+	0.2594	0.79235625		
+	0.2595	0.78940468		
+	0.2596	0.78453679		
+	0.2597	0.78408967		
+	0.2598	0.78153387		
+	0.2599	0.78387079		
+	0.26	0.7819896		
+	0.2601	0.80187232		
+	0.2602	0.80490027		
+	0.2603	0.80792366		
+	0.2604	0.82095711		
+	0.2605	0.83481995		
+	0.2606	0.83229288		
+	0.2607	0.84563478		
+	0.2608	0.84171115		
+	0.2609	0.8463178		
+	0.261	0.84185925		
+	0.2611	0.84408078		
+	0.2612	0.85900046		
+	0.2613	0.85644594		
+	0.2614	0.85756218		
+	0.2615	0.85865651		
+	0.2616	0.86183466		
+	0.2617	0.85956592		
+	0.2618	0.85816693		
+	0.2619	0.87322626		
+	0.262	0.8694028		
+	0.2621	0.86959671		
+	0.2622	0.86336508		
+	0.2623	0.87968287		
+	0.2624	0.88672678		
+	0.2625	0.8731308		
+	0.2626	0.88213808		
+	0.2627	0.88532821		
+	0.2628	0.88381088		
+	0.2629	0.88257173		
+	0.263	0.90430896		
+	0.2631	0.90146279		
+	0.2632	0.92431276		
+	0.2633	0.92123226		
+	0.2634	0.93996008		
+	0.2635	0.93428325		
+	0.2636	0.94776861		
+	0.2637	0.94060069		
+	0.2638	0.94765755		
+	0.2639	0.9430046		
+	0.264	0.94072185		
+	0.2641	0.93702254		
+	0.2642	0.9388631		
+	0.2643	0.92241801		
+	0.2644	0.92114195		
+	0.2645	0.93296787		
+	0.2646	0.92121053		
+	0.2647	0.91036156		
+	0.2648	0.91856823		
+	0.2649	0.9199857		
+	0.265	0.91427742		
+	0.2651	0.90031486		
+	0.2652	0.90692744		
+	0.2653	0.89081978		
+	0.2654	0.89465716		
+	0.2655	0.89067433		
+	0.2656	0.90046781		
+	0.2657	0.89067732		
+	0.2658	0.88912963		
+	0.2659	0.90476372		
+	0.266	0.9128219		
+	0.2661	0.92473553		
+	0.2662	0.93504579		
+	0.2663	0.93683206		
+	0.2664	0.94813086		
+	0.2665	0.95562131		
+	0.2666	0.95142451		
+	0.2667	0.95652327		
+	0.2668	0.93904954		
+	0.2669	0.93800592		
+	0.267	0.94369548		
+	0.2671	0.93459379		
+	0.2672	0.9420464		
+	0.2673	0.93596248		
+	0.2674	0.93264079		
+	0.2675	0.90918471		
+	0.2676	0.91681666		
+	0.2677	0.89504329		
+	0.2678	0.88539804		
+	0.2679	0.87523025		
+	0.268	0.86215261		
+	0.2681	0.85348932		
+	0.2682	0.84684501		
+	0.2683	0.84084793		
+	0.2684	0.84151239		
+	0.2685	0.81874538		
+	0.2686	0.82231758		
+	0.2687	0.81384333		
+	0.2688	0.83007587		
+	0.2689	0.82105655		
+	0.269	0.82433098		
+	0.2691	0.83476284		
+	0.2692	0.84499368		
+	0.2693	0.85372209		
+	0.2694	0.84690058		
+	0.2695	0.84809363		
+	0.2696	0.83341146		
+	0.2697	0.84101628		
+	0.2698	0.82674836		
+	0.2699	0.83197035		
+	0.27	0.82890616		
+	0.2701	0.81525374		
+	0.2702	0.81635778		
+	0.2703	0.82029498		
+	0.2704	0.8087204		
+	0.2705	0.8137556		
+	0.2706	0.79376008		
+	0.2707	0.79311703		
+	0.2708	0.7945514		
+	0.2709	0.78255973		
+	0.271	0.7925427		
+	0.2711	0.78717581		
+	0.2712	0.78289422		
+	0.2713	0.78339526		
+	0.2714	0.792792		
+	0.2715	0.77495866		
+	0.2716	0.77589758		
+	0.2717	0.79356371		
+	0.2718	0.78550515		
+	0.2719	0.79645231		
+	0.272	0.82525576		
+	0.2721	0.81784298		
+	0.2722	0.82314873		
+	0.2723	0.84197715		
+	0.2724	0.83284561		
+	0.2725	0.84121698		
+	0.2726	0.83002892		
+	0.2727	0.82827446		
+	0.2728	0.82635783		
+	0.2729	0.83453097		
+	0.273	0.82286527		
+	0.2731	0.82063166		
+	0.2732	0.81941986		
+	0.2733	0.81889727		
+	0.2734	0.81418293		
+	0.2735	0.79999537		
+	0.2736	0.79802668		
+	0.2737	0.79511271		
+	0.2738	0.79539132		
+	0.2739	0.79793956		
+	0.274	0.78796272		
+	0.2741	0.79002811		
+	0.2742	0.78375763		
+	0.2743	0.78968766		
+	0.2744	0.79145257		
+	0.2745	0.77834805		
+	0.2746	0.7927942		
+	0.2747	0.79790842		
+	0.2748	0.80325515		
+	0.2749	0.8257016		
+	0.275	0.82096579		
+	0.2751	0.83205729		
+	0.2752	0.84090911		
+	0.2753	0.83245495		
+	0.2754	0.83876055		
+	0.2755	0.83883359		
+	0.2756	0.83253004		
+	0.2757	0.83775375		
+	0.2758	0.82990504		
+	0.2759	0.82167769		
+	0.276	0.8201469		
+	0.2761	0.818528		
+	0.2762	0.81927092		
+	0.2763	0.80617081		
+	0.2764	0.81477678		
+	0.2765	0.8028795		
+	0.2766	0.80781637		
+	0.2767	0.79121276		
+	0.2768	0.79177822		
+	0.2769	0.79350508		
+	0.277	0.79789651		
+	0.2771	0.79450971		
+	0.2772	0.80519095		
+	0.2773	0.81018581		
+	0.2774	0.81281336		
+	0.2775	0.81166939		
+	0.2776	0.8221793		
+	0.2777	0.83342305		
+	0.2778	0.85074091		
+	0.2779	0.87694414		
+	0.278	0.892792		
+	0.2781	0.88379337		
+	0.2782	0.89642456		
+	0.2783	0.9159499		
+	0.2784	0.90211095		
+	0.2785	0.92395174		
+	0.2786	0.90976895		
+	0.2787	0.91963008		
+	0.2788	0.92301719		
+	0.2789	0.91324874		
+	0.279	0.92178794		
+	0.2791	0.91398424		
+	0.2792	0.90917251		
+	0.2793	0.90434279		
+	0.2794	0.8997756		
+	0.2795	0.90789042		
+	0.2796	0.90966166		
+	0.2797	0.90529491		
+	0.2798	0.90402705		
+	0.2799	0.89548286		
+	0.28	0.90373657		
+	0.2801	0.89804074		
+	0.2802	0.90409963		
+	0.2803	0.90349955		
+	0.2804	0.90098759		
+	0.2805	0.89482881		
+	0.2806	0.91738482		
+	0.2807	0.92627563		
+	0.2808	0.93080228		
+	0.2809	0.94853438		
+	0.281	0.95653865		
+	0.2811	0.94604329		
+	0.2812	0.95264816		
+	0.2813	0.95111192		
+	0.2814	0.94858448		
+	0.2815	0.94159646		
+	0.2816	0.94766895		
+	0.2817	0.94897222		
+	0.2818	0.94575772		
+	0.2819	0.93547727		
+	0.282	0.93937862		
+	0.2821	0.93572509		
+	0.2822	0.92597146		
+	0.2823	0.93067206		
+	0.2824	0.92268148		
+	0.2825	0.91318889		
+	0.2826	0.91372415		
+	0.2827	0.91754817		
+	0.2828	0.90997152		
+	0.2829	0.90385358		
+	0.283	0.90297668		
+	0.2831	0.89678093		
+	0.2832	0.91076361		
+	0.2833	0.89557966		
+	0.2834	0.91170736		
+	0.2835	0.9067882		
+	0.2836	0.9168436		
+	0.2837	0.93965109		
+	0.2838	0.93067793		
+	0.2839	0.93815635		
+	0.284	0.94579636		
+	0.2841	0.93522652		
+	0.2842	0.91235796		
+	0.2843	0.91168969		
+	0.2844	0.90436238		
+	0.2845	0.90501976		
+	0.2846	0.89721118		
+	0.2847	0.88187675		
+	0.2848	0.87999789		
+	0.2849	0.85882892		
+	0.285	0.85843291		
+	0.2851	0.85101061		
+	0.2852	0.84117691		
+	0.2853	0.82666352		
+	0.2854	0.82699373		
+	0.2855	0.82041691		
+	0.2856	0.80761311		
+	0.2857	0.80860208		
+	0.2858	0.80677708		
+	0.2859	0.80259283		
+	0.286	0.80073138		
+	0.2861	0.78474867		
+	0.2862	0.79745657		
+	0.2863	0.80184936		
+	0.2864	0.79657516		
+	0.2865	0.81230911		
+	0.2866	0.82571824		
+	0.2867	0.83017497		
+	0.2868	0.82909679		
+	0.2869	0.83862394		
+	0.287	0.84713779		
+	0.2871	0.83088579		
+	0.2872	0.83376978		
+	0.2873	0.83459909		
+	0.2874	0.84099339		
+	0.2875	0.83124719		
+	0.2876	0.82756673		
+	0.2877	0.83450199		
+	0.2878	0.81389228		
+	0.2879	0.82512766		
+	0.288	0.82200767		
+	0.2881	0.80457852		
+	0.2882	0.80062849		
+	0.2883	0.81163826		
+	0.2884	0.80905197		
+	0.2885	0.80691552		
+	0.2886	0.78660792		
+	0.2887	0.80256669		
+	0.2888	0.78429559		
+	0.2889	0.79472873		
+	0.289	0.79743248		
+	0.2891	0.78619023		
+	0.2892	0.79533616		
+	0.2893	0.79899841		
+	0.2894	0.80497786		
+	0.2895	0.82415552		
+	0.2896	0.83152885		
+	0.2897	0.83294838		
+	0.2898	0.83396862		
+	0.2899	0.84999864		
+	0.29	0.84615732		
+	0.2901	0.84338877		
+	0.2902	0.83891348		
+	0.2903	0.84255626		
+	0.2904	0.84524475		
+	0.2905	0.83721421		
+	0.2906	0.82304081		
+	0.2907	0.8175579		
+	0.2908	0.82715805		
+	0.2909	0.82761183		
+	0.291	0.81580169		
+	0.2911	0.80304413		
+	0.2912	0.8085169		
+	0.2913	0.81105826		
+	0.2914	0.80316069		
+	0.2915	0.79135534		
+	0.2916	0.79572166		
+	0.2917	0.79218463		
+	0.2918	0.79280454		
+	0.2919	0.79222862		
+	0.292	0.79724503		
+	0.2921	0.79999419		
+	0.2922	0.79742058		
+	0.2923	0.81466712		
+	0.2924	0.82630407		
+	0.2925	0.82495799		
+	0.2926	0.84349175		
+	0.2927	0.8501676		
+	0.2928	0.84378279		
+	0.2929	0.84379416		
+	0.293	0.84462484		
+	0.2931	0.8454787		
+	0.2932	0.85031388		
+	0.2933	0.83961711		
+	0.2934	0.85225698		
+	0.2935	0.84525497		
+	0.2936	0.84908526		
+	0.2937	0.83927584		
+	0.2938	0.84181046		
+	0.2939	0.83945356		
+	0.294	0.8408823		
+	0.2941	0.84705686		
+	0.2942	0.84628545		
+	0.2943	0.84702555		
+	0.2944	0.86175453		
+	0.2945	0.84891635		
+	0.2946	0.87084322		
+	0.2947	0.87494756		
+	0.2948	0.88096441		
+	0.2949	0.87952718		
+	0.295	0.87903072		
+	0.2951	0.8907409		
+	0.2952	0.89583814		
+	0.2953	0.91143107		
+	0.2954	0.92113029		
+	0.2955	0.93059513		
+	0.2956	0.93995269		
+	0.2957	0.94059086		
+	0.2958	0.95632891		
+	0.2959	0.93858385		
+	0.296	0.95684802		
+	0.2961	0.95242189		
+	0.2962	0.94403916		
+	0.2963	0.95296042		
+	0.2964	0.93271357		
+	0.2965	0.94352704		
+	0.2966	0.93259239		
+	0.2967	0.93544336		
+	0.2968	0.92341185		
+	0.2969	0.93361355		
+	0.297	0.9149895		
+	0.2971	0.92730445		
+	0.2972	0.90989808		
+	0.2973	0.91996233		
+	0.2974	0.90766787		
+	0.2975	0.91506046		
+	0.2976	0.91132266		
+	0.2977	0.90369034		
+	0.2978	0.91625617		
+	0.2979	0.91677839		
+	0.298	0.90942482		
+	0.2981	0.91873336		
+	0.2982	0.93088313		
+	0.2983	0.93687007		
+	0.2984	0.94294444		
+	0.2985	0.95855551		
+	0.2986	0.95049458		
+	0.2987	0.96699623		
+	0.2988	0.96586323		
+	0.2989	0.94990227		
+	0.299	0.95946155		
+	0.2991	0.94794699		
+	0.2992	0.95730616		
+	0.2993	0.94342684		
+	0.2994	0.95183839		
+	0.2995	0.95156505		
+	0.2996	0.94292027		
+	0.2997	0.93728985		
+	0.2998	0.93308427		
+	0.2999	0.92880866		
+	0.3	0.92016567		
+	0.3001	0.91983425		
+	0.3002	0.91430409		
+	0.3003	0.89634889		
+	0.3004	0.89281371		
+	0.3005	0.89400229		
+	0.3006	0.88428471		
+	0.3007	0.87529727		
+	0.3008	0.87048451		
+	0.3009	0.85161884		
+	0.301	0.86084975		
+	0.3011	0.8637884		
+	0.3012	0.86044866		
+	0.3013	0.87448058		
+	0.3014	0.86911048		
+	0.3015	0.88704558		
+	0.3016	0.88535894		
+	0.3017	0.86397846		
+	0.3018	0.8648591		
+	0.3019	0.86881008		
+	0.302	0.86731245		
+	0.3021	0.86271597		
+	0.3022	0.8441465		
+	0.3023	0.83712648		
+	0.3024	0.84173029		
+	0.3025	0.82601342		
+	0.3026	0.81907843		
+	0.3027	0.83245212		
+	0.3028	0.81194471		
+	0.3029	0.81843107		
+	0.303	0.81807641		
+	0.3031	0.79774931		
+	0.3032	0.81114041		
+	0.3033	0.80096211		
+	0.3034	0.79242482		
+	0.3035	0.80172634		
+	0.3036	0.79429535		
+	0.3037	0.79075744		
+	0.3038	0.79206199		
+	0.3039	0.80616788		
+	0.304	0.81054662		
+	0.3041	0.82594748		
+	0.3042	0.83369409		
+	0.3043	0.85221217		
+	0.3044	0.8505328		
+	0.3045	0.84038377		
+	0.3046	0.8449576		
+	0.3047	0.84037047		
+	0.3048	0.85442017		
+	0.3049	0.83600107		
+	0.305	0.84027827		
+	0.3051	0.84545327		
+	0.3052	0.83972981		
+	0.3053	0.83994475		
+	0.3054	0.82710436		
+	0.3055	0.83328753		
+	0.3056	0.82914304		
+	0.3057	0.81950412		
+	0.3058	0.82459884		
+	0.3059	0.8183193		
+	0.306	0.81642705		
+	0.3061	0.81609455		
+	0.3062	0.8034106		
+	0.3063	0.80999426		
+	0.3064	0.80827072		
+	0.3065	0.79646204		
+	0.3066	0.79703947		
+	0.3067	0.79564668		
+	0.3068	0.80075651		
+	0.3069	0.8049483		
+	0.307	0.81495756		
+	0.3071	0.8416478		
+	0.3072	0.85271153		
+	0.3073	0.84992567		
+	0.3074	0.86220697		
+	0.3075	0.85644592		
+	0.3076	0.853916		
+	0.3077	0.84962379		
+	0.3078	0.85036985		
+	0.3079	0.85135979		
+	0.308	0.84619478		
+	0.3081	0.84071211		
+	0.3082	0.84511514		
+	0.3083	0.83982277		
+	0.3084	0.83862228		
+	0.3085	0.81976609		
+	0.3086	0.82102327		
+	0.3087	0.82672604		
+	0.3088	0.81795341		
+	0.3089	0.80594656		
+	0.309	0.80950372		
+	0.3091	0.81290394		
+	0.3092	0.81688142		
+	0.3093	0.79825321		
+	0.3094	0.80888198		
+	0.3095	0.80121773		
+	0.3096	0.7998416		
+	0.3097	0.8116435		
+	0.3098	0.83389718		
+	0.3099	0.83981985		
+	0.31	0.86045513		
+	0.3101	0.87097085		
+	0.3102	0.87864421		
+	0.3103	0.88647598		
+	0.3104	0.88740303		
+	0.3105	0.89415319		
+	0.3106	0.90484777		
+	0.3107	0.89943404		
+	0.3108	0.90563666		
+	0.3109	0.91562149		
+	0.311	0.90396		
+	0.3111	0.91897281		
+	0.3112	0.91039598		
+	0.3113	0.9281798		
+	0.3114	0.92918647		
+	0.3115	0.92452631		
+	0.3116	0.90936348		
+	0.3117	0.91173548		
+	0.3118	0.92491533		
+	0.3119	0.90674157		
+	0.312	0.90952891		
+	0.3121	0.91128303		
+	0.3122	0.91193719		
+	0.3123	0.90172565		
+	0.3124	0.90999943		
+	0.3125	0.9006892		
+	0.3126	0.92067285		
+	0.3127	0.91512724		
+	0.3128	0.93125379		
+	0.3129	0.94071138		
+	0.313	0.9431663		
+	0.3131	0.95466482		
+	0.3132	0.97418174		
+	0.3133	0.96739626		
+	0.3134	0.96342044		
+	0.3135	0.96311778		
+	0.3136	0.95951352		
+	0.3137	0.96787777		
+	0.3138	0.95195808		
+	0.3139	0.95975961		
+	0.314	0.95755041		
+	0.3141	0.94322272		
+	0.3142	0.93880308		
+	0.3143	0.93877247		
+	0.3144	0.94048674		
+	0.3145	0.94381214		
+	0.3146	0.93532984		
+	0.3147	0.93555646		
+	0.3148	0.93388606		
+	0.3149	0.9297742		
+	0.315	0.92193775		
+	0.3151	0.91781165		
+	0.3152	0.91513474		
+	0.3153	0.91684516		
+	0.3154	0.91971475		
+	0.3155	0.91829655		
+	0.3156	0.92599083		
+	0.3157	0.93991361		
+	0.3158	0.94145088		
+	0.3159	0.9595627		
+	0.316	0.955809		
+	0.3161	0.97054076		
+	0.3162	0.97160443		
+	0.3163	0.97156159		
+	0.3164	0.97023456		
+	0.3165	0.96094009		
+	0.3166	0.95523643		
+	0.3167	0.95514358		
+	0.3168	0.94689175		
+	0.3169	0.92869156		
+	0.317	0.91019162		
+	0.3171	0.91386102		
+	0.3172	0.89540155		
+	0.3173	0.88769859		
+	0.3174	0.87174231		
+	0.3175	0.87946628		
+	0.3176	0.86771387		
+	0.3177	0.85700665		
+	0.3178	0.84702001		
+	0.3179	0.85127903		
+	0.318	0.83401001		
+	0.3181	0.83740878		
+	0.3182	0.82555093		
+	0.3183	0.82889795		
+	0.3184	0.82170611		
+	0.3185	0.83120655		
+	0.3186	0.82247077		
+	0.3187	0.84160628		
+	0.3188	0.85645434		
+	0.3189	0.85338531		
+	0.319	0.86828033		
+	0.3191	0.85460995		
+	0.3192	0.86875501		
+	0.3193	0.85689921		
+	0.3194	0.86401118		
+	0.3195	0.85342732		
+	0.3196	0.8556825		
+	0.3197	0.84838523		
+	0.3198	0.85466628		
+	0.3199	0.84554078		
+	0.32	0.8386524		
+	0.3201	0.84000015		
+	0.3202	0.82613088		
+	0.3203	0.83418108		
+	0.3204	0.83321053		
+	0.3205	0.82101524		
+	0.3206	0.81134608		
+	0.3207	0.81181662		
+	0.3208	0.80636293		
+	0.3209	0.81051123		
+	0.321	0.80870464		
+	0.3211	0.80738195		
+	0.3212	0.80660325		
+	0.3213	0.80792992		
+	0.3214	0.80631999		
+	0.3215	0.82323843		
+	0.3216	0.82664377		
+	0.3217	0.83228531		
+	0.3218	0.85728827		
+	0.3219	0.86646921		
+	0.322	0.85502822		
+	0.3221	0.85512894		
+	0.3222	0.86020684		
+	0.3223	0.86872356		
+	0.3224	0.84971983		
+	0.3225	0.85543353		
+	0.3226	0.84556485		
+	0.3227	0.8538901		
+	0.3228	0.85226567		
+	0.3229	0.83991186		
+	0.323	0.84133135		
+	0.3231	0.83520886		
+	0.3232	0.83352173		
+	0.3233	0.82265243		
+	0.3234	0.81939823		
+	0.3235	0.82060003		
+	0.3236	0.82815259		
+	0.3237	0.82040596		
+	0.3238	0.80973417		
+	0.3239	0.81363137		
+	0.324	0.81196287		
+	0.3241	0.81530156		
+	0.3242	0.80528142		
+	0.3243	0.81538106		
+	0.3244	0.82504776		
+	0.3245	0.82640954		
+	0.3246	0.84259723		
+	0.3247	0.85329547		
+	0.3248	0.85474047		
+	0.3249	0.86324442		
+	0.325	0.86676529		
+	0.3251	0.86703528		
+	0.3252	0.86405779		
+	0.3253	0.8709358		
+	0.3254	0.85945067		
+	0.3255	0.86184844		
+	0.3256	0.84863583		
+	0.3257	0.84718625		
+	0.3258	0.85884436		
+	0.3259	0.83885189		
+	0.326	0.84037373		
+	0.3261	0.85414604		
+	0.3262	0.83632147		
+	0.3263	0.83844414		
+	0.3264	0.84654636		
+	0.3265	0.84924484		
+	0.3266	0.83900038		
+	0.3267	0.84201855		
+	0.3268	0.8563054		
+	0.3269	0.8585149		
+	0.327	0.85369763		
+	0.3271	0.86850521		
+	0.3272	0.88155859		
+	0.3273	0.89195514		
+	0.3274	0.89519096		
+	0.3275	0.92177301		
+	0.3276	0.93573422		
+	0.3277	0.94993755		
+	0.3278	0.96216199		
+	0.3279	0.95226423		
+	0.328	0.97345587		
+	0.3281	0.9729453		
+	0.3282	0.96819623		
+	0.3283	0.96738765		
+	0.3284	0.96855961		
+	0.3285	0.96823129		
+	0.3286	0.96197813		
+	0.3287	0.95212198		
+	0.3288	0.94780214		
+	0.3289	0.94115236		
+	0.329	0.9434149		
+	0.3291	0.94841531		
+	0.3292	0.94120956		
+	0.3293	0.94021673		
+	0.3294	0.93204633		
+	0.3295	0.93354429		
+	0.3296	0.93573601		
+	0.3297	0.9303928		
+	0.3298	0.93122005		
+	0.3299	0.93181001		
+	0.33	0.93484194		
+	0.3301	0.93275543		
+	0.3302	0.93199697		
+	0.3303	0.93480814		
+	0.3304	0.95891729		
+	0.3305	0.96335319		
+	0.3306	0.97990131		
+	0.3307	0.97933592		
+	0.3308	0.97882755		
+	0.3309	0.97235312		
+	0.331	0.97843703		
+	0.3311	0.98182365		
+	0.3312	0.9811216		
+	0.3313	0.98337059		
+	0.3314	0.96885504		
+	0.3315	0.96063837		
+	0.3316	0.97480453		
+	0.3317	0.95872758		
+	0.3318	0.96535815		
+	0.3319	0.94981965		
+	0.332	0.95864287		
+	0.3321	0.94720485		
+	0.3322	0.94230278		
+	0.3323	0.94080157		
+	0.3324	0.93029169		
+	0.3325	0.93905601		
+	0.3326	0.94173478		
+	0.3327	0.93865387		
+	0.3328	0.92371179		
+	0.3329	0.92979359		
+	0.333	0.9173371		
+	0.3331	0.92426647		
+	0.3332	0.91728118		
+	0.3333	0.91493079		
+	0.3334	0.92826639		
+	0.3335	0.92654289		
+	0.3336	0.92675341		
+	0.3337	0.92275948		
+	0.3338	0.9167464		
+	0.3339	0.91624972		
+	0.334	0.91082243		
+	0.3341	0.89917367		
+	0.3342	0.89580365		
+	0.3343	0.89356374		
+	0.3344	0.87947218		
+	0.3345	0.88111194		
+	0.3346	0.86620078		
+	0.3347	0.86645989		
+	0.3348	0.86619545		
+	0.3349	0.85120709		
+	0.335	0.83895512		
+	0.3351	0.83622347		
+	0.3352	0.830987		
+	0.3353	0.83158672		
+	0.3354	0.81816432		
+	0.3355	0.8153074		
+	0.3356	0.82097716		
+	0.3357	0.82949969		
+	0.3358	0.82740445		
+	0.3359	0.82767384		
+	0.336	0.82832139		
+	0.3361	0.82672206		
+	0.3362	0.84293042		
+	0.3363	0.85592013		
+	0.3364	0.86234416		
+	0.3365	0.87014257		
+	0.3366	0.87193716		
+	0.3367	0.8750036		
+	0.3368	0.87093475		
+	0.3369	0.87466775		
+	0.337	0.85815268		
+	0.3371	0.86728453		
+	0.3372	0.8650782		
+	0.3373	0.86881246		
+	0.3374	0.85856477		
+	0.3375	0.84594721		
+	0.3376	0.86006477		
+	0.3377	0.85039513		
+	0.3378	0.83386323		
+	0.3379	0.84319408		
+	0.338	0.84294975		
+	0.3381	0.83026372		
+	0.3382	0.83862637		
+	0.3383	0.82463053		
+	0.3384	0.82235886		
+	0.3385	0.82118427		
+	0.3386	0.82931592		
+	0.3387	0.82813816		
+	0.3388	0.82100779		
+	0.3389	0.81893709		
+	0.339	0.83947159		
+	0.3391	0.84222743		
+	0.3392	0.84588039		
+	0.3393	0.86573628		
+	0.3394	0.86302393		
+	0.3395	0.87848835		
+	0.3396	0.88025083		
+	0.3397	0.86992153		
+	0.3398	0.86261527		
+	0.3399	0.87613194		
+	0.34	0.87247171		
+	0.3401	0.86063561		
+	0.3402	0.85917578		
+	0.3403	0.86113877		
+	0.3404	0.86229785		
+	0.3405	0.8492675		
+	0.3406	0.84897952		
+	0.3407	0.85195824		
+	0.3408	0.84416524		
+	0.3409	0.83115568		
+	0.341	0.82907864		
+	0.3411	0.82403473		
+	0.3412	0.82307269		
+	0.3413	0.83531679		
+	0.3414	0.82667905		
+	0.3415	0.82581059		
+	0.3416	0.82769086		
+	0.3417	0.81858685		
+	0.3418	0.82144037		
+	0.3419	0.82408488		
+	0.342	0.85047835		
+	0.3421	0.84831933		
+	0.3422	0.87095819		
+	0.3423	0.86846934		
+	0.3424	0.87527267		
+	0.3425	0.8863317		
+	0.3426	0.88527632		
+	0.3427	0.90006887		
+	0.3428	0.90287591		
+	0.3429	0.8910252		
+	0.343	0.9064131		
+	0.3431	0.91053157		
+	0.3432	0.91354995		
+	0.3433	0.91485075		
+	0.3434	0.91075348		
+	0.3435	0.9014043		
+	0.3436	0.90417264		
+	0.3437	0.91597297		
+	0.3438	0.91832332		
+	0.3439	0.92266871		
+	0.344	0.92030323		
+	0.3441	0.92156285		
+	0.3442	0.918051		
+	0.3443	0.9252367		
+	0.3444	0.91831034		
+	0.3445	0.92613437		
+	0.3446	0.92087602		
+	0.3447	0.93041767		
+	0.3448	0.92522953		
+	0.3449	0.94649352		
+	0.345	0.95245002		
+	0.3451	0.96207562		
+	0.3452	0.9806879		
+	0.3453	0.98940964		
+	0.3454	0.98069094		
+	0.3455	0.9811254		
+	0.3456	0.99412572		
+	0.3457	0.98701574		
+	0.3458	0.98124126		
+	0.3459	0.98961448		
+	0.346	0.97740114		
+	0.3461	0.97239532		
+	0.3462	0.96889237		
+	0.3463	0.97916158		
+	0.3464	0.97641977		
+	0.3465	0.9713518		
+	0.3466	0.95978632		
+	0.3467	0.96006388		
+	0.3468	0.96369449		
+	0.3469	0.95855792		
+	0.347	0.93971902		
+	0.3471	0.95180009		
+	0.3472	0.94001167		
+	0.3473	0.9506672		
+	0.3474	0.95063353		
+	0.3475	0.94665839		
+	0.3476	0.93931367		
+	0.3477	0.93683449		
+	0.3478	0.94804449		
+	0.3479	0.967031		
+	0.348	0.97853765		
+	0.3481	0.98900083		
+	0.3482	0.98574678		
+	0.3483	0.99864313		
+	0.3484	0.99860201		
+	0.3485	0.98684945		
+	0.3486	0.988476		
+	0.3487	0.98927985		
+	0.3488	0.9848301		
+	0.3489	0.98460835		
+	0.349	0.97499564		
+	0.3491	0.97963848		
+	0.3492	0.98114344		
+	0.3493	0.96886833		
+	0.3494	0.95533668		
+	0.3495	0.95268709		
+	0.3496	0.92980195		
+	0.3497	0.92134334		
+	0.3498	0.90554871		
+	0.3499	0.8999422		
+	0.35	0.89881916		
+	0.3501	0.89016567		
+	0.3502	0.87699453		
+	0.3503	0.87865729		
+	0.3504	0.87101844		
+	0.3505	0.85971642		
+	0.3506	0.85521363		
+	0.3507	0.85731682		
+	0.3508	0.87922905		
+	0.3509	0.88317523		
+	0.351	0.89683861		
+	0.3511	0.89217185		
+	0.3512	0.88498092		
+	0.3513	0.89326375		
+	0.3514	0.88144721		
+	0.3515	0.8925777		
+	0.3516	0.8807832		
+	0.3517	0.8860235		
+	0.3518	0.87280056		
+	0.3519	0.87071713		
+	0.352	0.87659748		
+	0.3521	0.86618253		
+	0.3522	0.87017395		
+	0.3523	0.84765343		
+	0.3524	0.84669421		
+	0.3525	0.8582931		
+	0.3526	0.84022423		
+	0.3527	0.83447967		
+	0.3528	0.84573689		
+	0.3529	0.83111063		
+	0.353	0.83554723		
+	0.3531	0.83351317		
+	0.3532	0.84052113		
+	0.3533	0.82851286		
+	0.3534	0.82681396		
+	0.3535	0.83559588		
+	0.3536	0.82874233		
+	0.3537	0.85335839		
+	0.3538	0.86408354		
+	0.3539	0.86872864		
+	0.354	0.88274444		
+	0.3541	0.88592008		
+	0.3542	0.87752782		
+	0.3543	0.87686513		
+	0.3544	0.87381618		
+	0.3545	0.88974722		
+	0.3546	0.88380595		
+	0.3547	0.87826049		
+	0.3548	0.8754434		
+	0.3549	0.86649309		
+	0.355	0.86103457		
+	0.3551	0.86902025		
+	0.3552	0.86407336		
+	0.3553	0.85547504		
+	0.3554	0.84756763		
+	0.3555	0.84463144		
+	0.3556	0.84517715		
+	0.3557	0.84213111		
+	0.3558	0.83519411		
+	0.3559	0.83428633		
+	0.356	0.83772678		
+	0.3561	0.84052021		
+	0.3562	0.83102188		
+	0.3563	0.84005685		
+	0.3564	0.84367075		
+	0.3565	0.83510343		
+	0.3566	0.84451289		
+	0.3567	0.85785172		
+	0.3568	0.87481311		
+	0.3569	0.87210559		
+	0.357	0.88459615		
+	0.3571	0.88393893		
+	0.3572	0.8899742		
+	0.3573	0.89438829		
+	0.3574	0.88760105		
+	0.3575	0.88427093		
+	0.3576	0.88316966		
+	0.3577	0.87412627		
+	0.3578	0.88354027		
+	0.3579	0.87319433		
+	0.358	0.86531027		
+	0.3581	0.86590954		
+	0.3582	0.86509898		
+	0.3583	0.85246552		
+	0.3584	0.86166679		
+	0.3585	0.85154204		
+	0.3586	0.85739647		
+	0.3587	0.84495676		
+	0.3588	0.85416106		
+	0.3589	0.85428458		
+	0.359	0.84887044		
+	0.3591	0.8568787		
+	0.3592	0.85081421		
+	0.3593	0.85817304		
+	0.3594	0.87725762		
+	0.3595	0.88045955		
+	0.3596	0.90549513		
+	0.3597	0.91918609		
+	0.3598	0.93754465		
+	0.3599	0.93297247		
+	0.36	0.95166344		
+	0.3601	0.96037824		
+	0.3602	0.96723036		
+	0.3603	0.96142818		
+	0.3604	0.96432121		
+	0.3605	0.97836775		
+	0.3606	0.97357568		
+	0.3607	0.97493472		
+	0.3608	0.97758262		
+	0.3609	0.98058606		
+	0.361	0.97735178		
+	0.3611	0.96934438		
+	0.3612	0.95845561		
+	0.3613	0.96847303		
+	0.3614	0.9594437		
+	0.3615	0.94381184		
+	0.3616	0.94627534		
+	0.3617	0.95190002		
+	0.3618	0.95847115		
+	0.3619	0.94351358		
+	0.362	0.94530356		
+	0.3621	0.94598294		
+	0.3622	0.94160277		
+	0.3623	0.94986435		
+	0.3624	0.96347364		
+	0.3625	0.96764694		
+	0.3626	0.9749259		
+	0.3627	0.98227446		
+	0.3628	0.99654798		
+	0.3629	1.0059446		
+	0.363	1.0087009		
+	0.3631	1.0095013		
+	0.3632	1.0090566		
+	0.3633	1.0040673		
+	0.3634	0.99912915		
+	0.3635	1.0015887		
+	0.3636	0.98427422		
+	0.3637	0.99724423		
+	0.3638	0.99529258		
+	0.3639	0.97494902		
+	0.364	0.97396322		
+	0.3641	0.97596954		
+	0.3642	0.97727265		
+	0.3643	0.95908943		
+	0.3644	0.97424955		
+	0.3645	0.95248524		
+	0.3646	0.9503848		
+	0.3647	0.9516958		
+	0.3648	0.96105548		
+	0.3649	0.95703273		
+	0.365	0.96025778		
+	0.3651	0.94699256		
+	0.3652	0.95390215		
+	0.3653	0.95308873		
+	0.3654	0.95700633		
+	0.3655	0.97301863		
+	0.3656	0.9861027		
+	0.3657	0.98859237		
+	0.3658	0.99361848		
+	0.3659	0.97504303		
+	0.366	0.96555811		
+	0.3661	0.97213684		
+	0.3662	0.95558913		
+	0.3663	0.94960052		
+	0.3664	0.9374318		
+	0.3665	0.92597769		
+	0.3666	0.9310983		
+	0.3667	0.92415017		
+	0.3668	0.90684232		
+	0.3669	0.89690372		
+	0.367	0.89564304		
+	0.3671	0.88568423		
+	0.3672	0.87491506		
+	0.3673	0.87900508		
+	0.3674	0.86293667		
+	0.3675	0.87120823		
+	0.3676	0.8535451		
+	0.3677	0.84788502		
+	0.3678	0.85470173		
+	0.3679	0.84078379		
+	0.368	0.84343099		
+	0.3681	0.83515379		
+	0.3682	0.84698342		
+	0.3683	0.85637299		
+	0.3684	0.87010744		
+	0.3685	0.86760727		
+	0.3686	0.89097577		
+	0.3687	0.89530255		
+	0.3688	0.89331018		
+	0.3689	0.89192858		
+	0.369	0.882126		
+	0.3691	0.89160541		
+	0.3692	0.88771301		
+	0.3693	0.88365241		
+	0.3694	0.88691055		
+	0.3695	0.87177704		
+	0.3696	0.86843488		
+	0.3697	0.87099499		
+	0.3698	0.86789525		
+	0.3699	0.87323119		
+	0.37	0.85555238		
+	0.3701	0.85317335		
+	0.3702	0.85277639		
+	0.3703	0.85288487		
+	0.3704	0.85367155		
+	0.3705	0.84024991		
+	0.3706	0.85467515		
+	0.3707	0.84246166		
+	0.3708	0.8337672		
+	0.3709	0.84868966		
+	0.371	0.83947796		
+	0.3711	0.85331266		
+	0.3712	0.84528157		
+	0.3713	0.85625386		
+	0.3714	0.87693477		
+	0.3715	0.88737426		
+	0.3716	0.89917459		
+	0.3717	0.89141651		
+	0.3718	0.88842991		
+	0.3719	0.902248		
+	0.372	0.88627799		
+	0.3721	0.89921869		
+	0.3722	0.880001		
+	0.3723	0.88475364		
+	0.3724	0.89002861		
+	0.3725	0.88644592		
+	0.3726	0.8672011		
+	0.3727	0.86575679		
+	0.3728	0.87094046		
+	0.3729	0.86293883		
+	0.373	0.86938665		
+	0.3731	0.86680827		
+	0.3732	0.85900747		
+	0.3733	0.84928955		
+	0.3734	0.84088048		
+	0.3735	0.85010026		
+	0.3736	0.84160724		
+	0.3737	0.83897958		
+	0.3738	0.83468689		
+	0.3739	0.84533784		
+	0.374	0.85703113		
+	0.3741	0.84737629		
+	0.3742	0.87301607		
+	0.3743	0.87309999		
+	0.3744	0.89075445		
+	0.3745	0.88516555		
+	0.3746	0.89746284		
+	0.3747	0.90344124		
+	0.3748	0.90099266		
+	0.3749	0.89925821		
+	0.375	0.88795021		
+	0.3751	0.90403708		
+	0.3752	0.90774488		
+	0.3753	0.8938944		
+	0.3754	0.89013604		
+	0.3755	0.90336545		
+	0.3756	0.89902878		
+	0.3757	0.90339949		
+	0.3758	0.91060338		
+	0.3759	0.90749444		
+	0.376	0.89675575		
+	0.3761	0.91406259		
+	0.3762	0.90685809		
+	0.3763	0.91878699		
+	0.3764	0.91089717		
+	0.3765	0.91436821		
+	0.3766	0.92742872		
+	0.3767	0.93083375		
+	0.3768	0.93751497		
+	0.3769	0.93010463		
+	0.377	0.9441855		
+	0.3771	0.95832331		
+	0.3772	0.97861624		
+	0.3773	0.9914035		
+	0.3774	0.99241995		
+	0.3775	0.99034515		
+	0.3776	0.9978277		
+	0.3777	0.99623055		
+	0.3778	1.0040743		
+	0.3779	0.99324416		
+	0.378	0.98829543		
+	0.3781	0.99737377		
+	0.3782	0.99657238		
+	0.3783	0.98737657		
+	0.3784	0.99853813		
+	0.3785	0.98380859		
+	0.3786	0.99300503		
+	0.3787	0.98606348		
+	0.3788	0.97617318		
+	0.3789	0.97807819		
+	0.379	0.96704491		
+	0.3791	0.97362074		
+	0.3792	0.97097601		
+	0.3793	0.95961769		
+	0.3794	0.95620682		
+	0.3795	0.95588203		
+	0.3796	0.96250303		
+	0.3797	0.95198098		
+	0.3798	0.96060604		
+	0.3799	0.97517427		
+	0.38	0.98232455		
+	0.3801	0.99280745		
+	0.3802	1.0033797		
+	0.3803	0.99825391		
+	0.3804	1.009656		
+	0.3805	1.0205142		
+	0.3806	1.0171518		
+	0.3807	1.0099893		
+	0.3808	1.0115071		
+	0.3809	1.0004694		
+	0.381	1.0112798		
+	0.3811	1.0145105		
+	0.3812	1.0017034		
+	0.3813	0.99506548		
+	0.3814	0.98569304		
+	0.3815	0.98230158		
+	0.3816	0.98236142		
+	0.3817	0.98275791		
+	0.3818	0.9764875		
+	0.3819	0.98020082		
+	0.382	0.96506139		
+	0.3821	0.95224902		
+	0.3822	0.96082524		
+	0.3823	0.93762295		
+	0.3824	0.92656515		
+	0.3825	0.93125043		
+	0.3826	0.91143542		
+	0.3827	0.90477112		
+	0.3828	0.91872997		
+	0.3829	0.91911956		
+	0.383	0.92010303		
+	0.3831	0.92028311		
+	0.3832	0.91984934		
+	0.3833	0.93809743		
+	0.3834	0.92060255		
+	0.3835	0.93175991		
+	0.3836	0.9182615		
+	0.3837	0.91951856		
+	0.3838	0.90714985		
+	0.3839	0.9032741		
+	0.384	0.91356833		
+	0.3841	0.89466167		
+	0.3842	0.89774882		
+	0.3843	0.88882507		
+	0.3844	0.89239079		
+	0.3845	0.88426727		
+	0.3846	0.88202122		
+	0.3847	0.86584613		
+	0.3848	0.86619421		
+	0.3849	0.85738303		
+	0.385	0.85945762		
+	0.3851	0.84865755		
+	0.3852	0.85608502		
+	0.3853	0.84390307		
+	0.3854	0.8428851		
+	0.3855	0.8431947		
+	0.3856	0.8542393		
+	0.3857	0.85712122		
+	0.3858	0.8523204		
+	0.3859	0.86140202		
+	0.386	0.86914305		
+	0.3861	0.89189011		
+	0.3862	0.89666109		
+	0.3863	0.89329456		
+	0.3864	0.89600004		
+	0.3865	0.89788389		
+	0.3866	0.90331851		
+	0.3867	0.89122706		
+	0.3868	0.89959866		
+	0.3869	0.90091616		
+	0.387	0.897701		
+	0.3871	0.87778064		
+	0.3872	0.87852032		
+	0.3873	0.88880285		
+	0.3874	0.86898541		
+	0.3875	0.87362238		
+	0.3876	0.87044851		
+	0.3877	0.85745601		
+	0.3878	0.86646033		
+	0.3879	0.85707666		
+	0.388	0.84805206		
+	0.3881	0.85483309		
+	0.3882	0.85844106		
+	0.3883	0.85531011		
+	0.3884	0.85795848		
+	0.3885	0.85153454		
+	0.3886	0.86101923		
+	0.3887	0.85542729		
+	0.3888	0.86244123		
+	0.3889	0.88052232		
+	0.389	0.89029871		
+	0.3891	0.90501886		
+	0.3892	0.9001147		
+	0.3893	0.90615377		
+	0.3894	0.8971847		
+	0.3895	0.9102549		
+	0.3896	0.90738701		
+	0.3897	0.89527141		
+	0.3898	0.90311578		
+	0.3899	0.89336302		
+	0.39	0.89007003		
+	0.3901	0.89599312		
+	0.3902	0.88899049		
+	0.3903	0.88225895		
+	0.3904	0.88242044		
+	0.3905	0.86763131		
+	0.3906	0.86339926		
+	0.3907	0.86733633		
+	0.3908	0.86839955		
+	0.3909	0.85098724		
+	0.391	0.84949446		
+	0.3911	0.86242402		
+	0.3912	0.86346119		
+	0.3913	0.85471415		
+	0.3914	0.85676005		
+	0.3915	0.85087579		
+	0.3916	0.87550994		
+	0.3917	0.8724705		
+	0.3918	0.90090121		
+	0.3919	0.91416137		
+	0.392	0.92458819		
+	0.3921	0.92978401		
+	0.3922	0.93995859		
+	0.3923	0.94972379		
+	0.3924	0.94955302		
+	0.3925	0.9430884		
+	0.3926	0.96324202		
+	0.3927	0.96485017		
+	0.3928	0.95353115		
+	0.3929	0.97390608		
+	0.393	0.97382245		
+	0.3931	0.97524171		
+	0.3932	0.96760128		
+	0.3933	0.96759081		
+	0.3934	0.97477551		
+	0.3935	0.96321882		
+	0.3936	0.9657004		
+	0.3937	0.9576082		
+	0.3938	0.96737087		
+	0.3939	0.96232577		
+	0.394	0.96021572		
+	0.3941	0.96682183		
+	0.3942	0.95018162		
+	0.3943	0.94844025		
+	0.3944	0.95574118		
+	0.3945	0.95664374		
+	0.3946	0.9740521		
+	0.3947	0.98989163		
+	0.3948	0.98561413		
+	0.3949	0.99404493		
+	0.395	1.0154628		
+	0.3951	1.0169458		
+	0.3952	1.008733		
+	0.3953	1.0070296		
+	0.3954	1.0224084		
+	0.3955	1.0139589		
+	0.3956	1.0137135		
+	0.3957	1.0089896		
+	0.3958	1.0059751		
+	0.3959	1.008558		
+	0.396	0.99710642		
+	0.3961	0.98949479		
+	0.3962	0.99115762		
+	0.3963	0.98523573		
+	0.3964	0.98069029		
+	0.3965	0.98109304		
+	0.3966	0.97724064		
+	0.3967	0.97001541		
+	0.3968	0.97689206		
+	0.3969	0.96535605		
+	0.397	0.96877816		
+	0.3971	0.96281228		
+	0.3972	0.96302017		
+	0.3973	0.9625999		
+	0.3974	0.96134005		
+	0.3975	0.97713691		
+	0.3976	0.97899777		
+	0.3977	0.99447513		
+	0.3978	0.99788023		
+	0.3979	1.0211598		
+	0.398	1.0228949		
+	0.3981	1.0246265		
+	0.3982	1.0233359		
+	0.3983	1.0192839		
+	0.3984	1.0042639		
+	0.3985	1.0062633		
+	0.3986	1.0013763		
+	0.3987	0.99220769		
+	0.3988	0.97150461		
+	0.3989	0.96305191		
+	0.399	0.95092972		
+	0.3991	0.94495558		
+	0.3992	0.93787191		
+	0.3993	0.92033074		
+	0.3994	0.92473751		
+	0.3995	0.90887584		
+	0.3996	0.90323568		
+	0.3997	0.89722273		
+	0.3998	0.89197928		
+	0.3999	0.89251602		
+	0.4	0.88403277		
+	0.4001	0.86471682		
+	0.4002	0.86847709		
+	0.4003	0.8637073		
+	0.4004	0.87951196		
+	0.4005	0.87718727		
+	0.4006	0.89078171		
+	0.4007	0.88753308		
+	0.4008	0.90574306		
+	0.4009	0.90005127		
+	0.401	0.9028892		
+	0.4011	0.90701361		
+	0.4012	0.89677537		
+	0.4013	0.89804449		
+	0.4014	0.90641288		
+	0.4015	0.90484671		
+	0.4016	0.88992295		
+	0.4017	0.88475322		
+	0.4018	0.88195561		
+	0.4019	0.88871341		
+	0.402	0.88022034		
+	0.4021	0.86694307		
+	0.4022	0.8744806		
+	0.4023	0.87008593		
+	0.4024	0.87132169		
+	0.4025	0.87102049		
+	0.4026	0.85943783		
+	0.4027	0.85117018		
+	0.4028	0.85141118		
+	0.4029	0.86414076		
+	0.403	0.85384671		
+	0.4031	0.84828099		
+	0.4032	0.84836322		
+	0.4033	0.84980511		
+	0.4034	0.8689493		
+	0.4035	0.87362447		
+	0.4036	0.88168894		
+	0.4037	0.88930698		
+	0.4038	0.89687245		
+	0.4039	0.90573011		
+	0.404	0.91194822		
+	0.4041	0.89437611		
+	0.4042	0.89469985		
+	0.4043	0.90188273		
+	0.4044	0.89668778		
+	0.4045	0.90084639		
+	0.4046	0.89397888		
+	0.4047	0.89499901		
+	0.4048	0.89129002		
+	0.4049	0.88327915		
+	0.405	0.87088941		
+	0.4051	0.87992762		
+	0.4052	0.86183613		
+	0.4053	0.86857708		
+	0.4054	0.86027731		
+	0.4055	0.85476048		
+	0.4056	0.85440122		
+	0.4057	0.85751303		
+	0.4058	0.85866191		
+	0.4059	0.84732903		
+	0.406	0.84901447		
+	0.4061	0.84886346		
+	0.4062	0.85855079		
+	0.4063	0.85906022		
+	0.4064	0.88205823		
+	0.4065	0.89175276		
+	0.4066	0.90301458		
+	0.4067	0.8988075		
+	0.4068	0.90276257		
+	0.4069	0.91529374		
+	0.407	0.90876475		
+	0.4071	0.91239903		
+	0.4072	0.90819752		
+	0.4073	0.90619027		
+	0.4074	0.89676616		
+	0.4075	0.88747535		
+	0.4076	0.90188779		
+	0.4077	0.88194711		
+	0.4078	0.88009812		
+	0.4079	0.89626		
+	0.408	0.88547845		
+	0.4081	0.89358507		
+	0.4082	0.87784301		
+	0.4083	0.89604995		
+	0.4084	0.89482742		
+	0.4085	0.89643895		
+	0.4086	0.88983028		
+	0.4087	0.90025077		
+	0.4088	0.89439396		
+	0.4089	0.91372234		
+	0.409	0.91716645		
+	0.4091	0.91415025		
+	0.4092	0.93671608		
+	0.4093	0.95803492		
+	0.4094	0.96548487		
+	0.4095	0.98152502		
+	0.4096	0.98748957		
+	0.4097	1.0023144		
+	0.4098	0.99335857		
+	0.4099	1.0055595		
+	0.41	1.0080008		
+	0.4101	0.99906851		
+	0.4102	1.008939		
+	0.4103	0.99531488		
+	0.4104	1.0017793		
+	0.4105	0.99061605		
+	0.4106	0.99422149		
+	0.4107	0.98099071		
+	0.4108	0.99354366		
+	0.4109	0.97387043		
+	0.411	0.97109604		
+	0.4111	0.98391866		
+	0.4112	0.96645074		
+	0.4113	0.96766092		
+	0.4114	0.96241146		
+	0.4115	0.97323147		
+	0.4116	0.96326004		
+	0.4117	0.96444852		
+	0.4118	0.96199157		
+	0.4119	0.96594576		
+	0.412	0.97755079		
+	0.4121	0.97342294		
+	0.4122	0.98449217		
+	0.4123	0.9945862		
+	0.4124	1.0123248		
+	0.4125	1.0181802		
+	0.4126	1.0162234		
+	0.4127	1.0195914		
+	0.4128	1.0169043		
+	0.4129	1.017646		
+	0.413	1.0202669		
+	0.4131	1.0141133		
+	0.4132	1.0089409		
+	0.4133	1.0011175		
+	0.4134	1.0166907		
+	0.4135	1.0045484		
+	0.4136	1.0087534		
+	0.4137	0.98963415		
+	0.4138	0.98709348		
+	0.4139	0.99236418		
+	0.414	0.98370449		
+	0.4141	0.98720196		
+	0.4142	0.98311218		
+	0.4143	0.98552318		
+	0.4144	0.97420112		
+	0.4145	0.97682053		
+	0.4146	0.96338115		
+	0.4147	0.9585442		
+	0.4148	0.95813911		
+	0.4149	0.95949826		
+	0.415	0.96591661		
+	0.4151	0.96708158		
+	0.4152	0.95678148		
+	0.4153	0.95722357		
+	0.4154	0.97134498		
+	0.4155	0.97257062		
+	0.4156	0.96490203		
+	0.4157	0.95426688		
+	0.4158	0.96114961		
+	0.4159	0.94576524		
+	0.416	0.93031041		
+	0.4161	0.92427976		
+	0.4162	0.9309197		
+	0.4163	0.92783058		
+	0.4164	0.91714505		
+	0.4165	0.90129465		
+	0.4166	0.90410827		
+	0.4167	0.89028001		
+	0.4168	0.89264001		
+	0.4169	0.88185012		
+	0.417	0.86665202		
+	0.4171	0.87350596		
+	0.4172	0.86042619		
+	0.4173	0.86440689		
+	0.4174	0.85200043		
+	0.4175	0.86131663		
+	0.4176	0.86000369		
+	0.4177	0.84641035		
+	0.4178	0.86362966		
+	0.4179	0.85124343		
+	0.418	0.86267919		
+	0.4181	0.87414967		
+	0.4182	0.87974233		
+	0.4183	0.88734811		
+	0.4184	0.89402283		
+	0.4185	0.91326339		
+	0.4186	0.91396873		
+	0.4187	0.9088738		
+	0.4188	0.89589394		
+	0.4189	0.8931819		
+	0.419	0.90306265		
+	0.4191	0.89223547		
+	0.4192	0.89447733		
+	0.4193	0.88218963		
+	0.4194	0.88885826		
+	0.4195	0.87874459		
+	0.4196	0.87911634		
+	0.4197	0.87205398		
+	0.4198	0.86442762		
+	0.4199	0.86621484		
+	0.42	0.8556625		
+	0.4201	0.85870981		
+	0.4202	0.87013259		
+	0.4203	0.8563758		
+	0.4204	0.84899299		
+	0.4205	0.8484785		
+	0.4206	0.85387512		
+	0.4207	0.85249921		
+	0.4208	0.85199258		
+	0.4209	0.87291593		
+	0.421	0.88164154		
+	0.4211	0.89452604		
+	0.4212	0.89514897		
+	0.4213	0.90771959		
+	0.4214	0.89924174		
+	0.4215	0.9128287		
+	0.4216	0.91138868		
+	0.4217	0.90265723		
+	0.4218	0.90598565		
+	0.4219	0.89258282		
+	0.422	0.89695536		
+	0.4221	0.89173987		
+	0.4222	0.89868548		
+	0.4223	0.88022123		
+	0.4224	0.8878406		
+	0.4225	0.89193959		
+	0.4226	0.87398524		
+	0.4227	0.8710442		
+	0.4228	0.8621353		
+	0.4229	0.86475374		
+	0.423	0.86565301		
+	0.4231	0.87219975		
+	0.4232	0.85161821		
+	0.4233	0.85679861		
+	0.4234	0.8472178		
+	0.4235	0.85381699		
+	0.4236	0.85053511		
+	0.4237	0.86218532		
+	0.4238	0.85983256		
+	0.4239	0.87874616		
+	0.424	0.89316338		
+	0.4241	0.88755369		
+	0.4242	0.91419345		
+	0.4243	0.92120372		
+	0.4244	0.92355483		
+	0.4245	0.92500894		
+	0.4246	0.91505825		
+	0.4247	0.93200164		
+	0.4248	0.9298734		
+	0.4249	0.93243675		
+	0.425	0.93329289		
+	0.4251	0.93365649		
+	0.4252	0.93262957		
+	0.4253	0.94281171		
+	0.4254	0.94151595		
+	0.4255	0.93340351		
+	0.4256	0.94253499		
+	0.4257	0.94845265		
+	0.4258	0.94124248		
+	0.4259	0.95261857		
+	0.426	0.94291645		
+	0.4261	0.9503681		
+	0.4262	0.94569986		
+	0.4263	0.95831578		
+	0.4264	0.94630041		
+	0.4265	0.95071193		
+	0.4266	0.96331676		
+	0.4267	0.96378215		
+	0.4268	0.97063351		
+	0.4269	0.97583436		
+	0.427	0.99724126		
+	0.4271	0.99635861		
+	0.4272	1.0085324		
+	0.4273	1.0085477		
+	0.4274	1.0179888		
+	0.4275	1.0181131		
+	0.4276	1.0047159		
+	0.4277	1.0116317		
+	0.4278	1.0177376		
+	0.4279	1.0066632		
+	0.428	0.99485114		
+	0.4281	1.0057158		
+	0.4282	1.0043851		
+	0.4283	0.98935431		
+	0.4284	0.99689924		
+	0.4285	0.98680798		
+	0.4286	0.98120279		
+	0.4287	0.9776451		
+	0.4288	0.97802194		
+	0.4289	0.97139058		
+	0.429	0.97198554		
+	0.4291	0.97268988		
+	0.4292	0.97531103		
+	0.4293	0.96087123		
+	0.4294	0.97424912		
+	0.4295	0.95985843		
+	0.4296	0.96947512		
+	0.4297	0.98988435		
+	0.4298	0.99299751		
+	0.4299	1.0111377		
+	0.43	1.0047204		
+	0.4301	1.0146167		
+	0.4302	1.0132594		
+	0.4303	1.0161119		
+	0.4304	1.0182383		
+	0.4305	1.0157891		
+	0.4306	1.0227108		
+	0.4307	1.0173321		
+	0.4308	1.0111715		
+	0.4309	1.0160993		
+	0.431	1.0036656		
+	0.4311	0.99786963		
+	0.4312	0.98661519		
+	0.4313	0.98180798		
+	0.4314	0.97866488		
+	0.4315	0.95569983		
+	0.4316	0.95039388		
+	0.4317	0.93783105		
+	0.4318	0.92263018		
+	0.4319	0.91748222		
+	0.432	0.90758202		
+	0.4321	0.9051601		
+	0.4322	0.89349593		
+	0.4323	0.90409757		
+	0.4324	0.89569579		
+	0.4325	0.88954347		
+	0.4326	0.89396205		
+	0.4327	0.90646346		
+	0.4328	0.90592998		
+	0.4329	0.91335272		
+	0.433	0.91905929		
+	0.4331	0.91347255		
+	0.4332	0.92369232		
+	0.4333	0.90366748		
+	0.4334	0.91630135		
+	0.4335	0.91233191		
+	0.4336	0.90139449		
+	0.4337	0.89909194		
+	0.4338	0.88865272		
+	0.4339	0.88287312		
+	0.434	0.88147287		
+	0.4341	0.88928467		
+	0.4342	0.88200355		
+	0.4343	0.88195282		
+	0.4344	0.86580569		
+	0.4345	0.86225101		
+	0.4346	0.85864864		
+	0.4347	0.86434826		
+	0.4348	0.85518339		
+	0.4349	0.85377975		
+	0.435	0.84833161		
+	0.4351	0.86069798		
+	0.4352	0.85599019		
+	0.4353	0.85178773		
+	0.4354	0.85078367		
+	0.4355	0.8562266		
+	0.4356	0.86968413		
+	0.4357	0.8820472		
+	0.4358	0.89146864		
+	0.4359	0.9000352		
+	0.436	0.89554565		
+	0.4361	0.90316908		
+	0.4362	0.90262978		
+	0.4363	0.89990404		
+	0.4364	0.9051771		
+	0.4365	0.90731408		
+	0.4366	0.89961095		
+	0.4367	0.89698296		
+	0.4368	0.88401282		
+	0.4369	0.88752295		
+	0.437	0.88453127		
+	0.4371	0.87815401		
+	0.4372	0.88518083		
+	0.4373	0.86472251		
+	0.4374	0.87375063		
+	0.4375	0.86866431		
+	0.4376	0.85355949		
+	0.4377	0.8489739		
+	0.4378	0.85999023		
+	0.4379	0.84810711		
+	0.438	0.85540745		
+	0.4381	0.85299256		
+	0.4382	0.85126198		
+	0.4383	0.85852369		
+	0.4384	0.86492639		
+	0.4385	0.86610134		
+	0.4386	0.86930049		
+	0.4387	0.89446039		
+	0.4388	0.90152109		
+	0.4389	0.90637637		
+	0.439	0.9045957		
+	0.4391	0.90149741		
+	0.4392	0.90386976		
+	0.4393	0.90716204		
+	0.4394	0.9084793		
+	0.4395	0.90629463		
+	0.4396	0.88904871		
+	0.4397	0.89780468		
+	0.4398	0.89626238		
+	0.4399	0.88253208		
+	0.44	0.8817951		
+	0.4401	0.86851726		
+	0.4402	0.87661586		
+	0.4403	0.87791722		
+	0.4404	0.86933608		
+	0.4405	0.87120335		
+	0.4406	0.87246528		
+	0.4407	0.87005739		
+	0.4408	0.87071951		
+	0.4409	0.8737297		
+	0.441	0.86261856		
+	0.4411	0.87019336		
+	0.4412	0.87729866		
+	0.4413	0.89727278		
+	0.4414	0.8922964		
+	0.4415	0.91983746		
+	0.4416	0.93785158		
+	0.4417	0.94433043		
+	0.4418	0.9667478		
+	0.4419	0.97047986		
+	0.442	0.96531497		
+	0.4421	0.98505131		
+	0.4422	0.98872847		
+	0.4423	0.98135737		
+	0.4424	0.99163499		
+	0.4425	0.98448622		
+	0.4426	0.99388329		
+	0.4427	0.98920636		
+	0.4428	0.97619454		
+	0.4429	0.9880168		
+	0.443	0.98050484		
+	0.4431	0.96675057		
+	0.4432	0.96702007		
+	0.4433	0.96531631		
+	0.4434	0.96437336		
+	0.4435	0.95875874		
+	0.4436	0.97078717		
+	0.4437	0.95321247		
+	0.4438	0.95093162		
+	0.4439	0.9682274		
+	0.444	0.95220372		
+	0.4441	0.96668509		
+	0.4442	0.9661411		
+	0.4443	0.9810455		
+	0.4444	0.97245882		
+	0.4445	0.99456855		
+	0.4446	0.9964304		
+	0.4447	1.0024236		
+	0.4448	1.0132057		
+	0.4449	1.0072665		
+	0.445	1.0151557		
+	0.4451	1.0171386		
+	0.4452	1.0051989		
+	0.4453	1.007585		
+	0.4454	1.0128061		
+	0.4455	1.0043287		
+	0.4456	1.0061706		
+	0.4457	1.0036799		
+	0.4458	0.99304904		
+	0.4459	0.99283838		
+	0.446	0.99213716		
+	0.4461	0.98943891		
+	0.4462	0.97056618		
+	0.4463	0.9757836		
+	0.4464	0.96517213		
+	0.4465	0.96874283		
+	0.4466	0.96178308		
+	0.4467	0.97108019		
+	0.4468	0.96161902		
+	0.4469	0.97140181		
+	0.447	0.96687022		
+	0.4471	0.96009125		
+	0.4472	0.97669141		
+	0.4473	0.98299304		
+	0.4474	0.99344622		
+	0.4475	1.0016052		
+	0.4476	1.0008819		
+	0.4477	0.99757826		
+	0.4478	0.98925169		
+	0.4479	0.98074134		
+	0.448	0.98245332		
+	0.4481	0.97601769		
+	0.4482	0.95745464		
+	0.4483	0.95441237		
+	0.4484	0.94398014		
+	0.4485	0.94412313		
+	0.4486	0.9365009		
+	0.4487	0.91506554		
+	0.4488	0.91917089		
+	0.4489	0.89496111		
+	0.449	0.89602043		
+	0.4491	0.89398484		
+	0.4492	0.88006292		
+	0.4493	0.87268341		
+	0.4494	0.87932373		
+	0.4495	0.8727868		
+	0.4496	0.86854085		
+	0.4497	0.86167644		
+	0.4498	0.86167563		
+	0.4499	0.84777898		
+	0.45	0.86167563		
+	0.4501	0.85003242		
+	0.4502	0.8743317		
+	0.4503	0.8688096		
+	0.4504	0.87784683		
+	0.4505	0.89002637		
+	0.4506	0.90001168		
+	0.4507	0.89416032		
+	0.4508	0.90515944		
+	0.4509	0.90261909		
+	0.451	0.88914774		
+	0.4511	0.89067291		
+	0.4512	0.88982202		
+	0.4513	0.88866055		
+	0.4514	0.88786546		
+	0.4515	0.87370911		
+	0.4516	0.88472368		
+	0.4517	0.87975316		
+	0.4518	0.86384953		
+	0.4519	0.87262132		
+	0.452	0.86320019		
+	0.4521	0.85767371		
+	0.4522	0.84804775		
+	0.4523	0.84674305		
+	0.4524	0.849995		
+	0.4525	0.83988514		
+	0.4526	0.84705168		
+	0.4527	0.85097419		
+	0.4528	0.84909949		
+	0.4529	0.84028385		
+	0.453	0.84234514		
+	0.4531	0.85163702		
+	0.4532	0.87674074		
+	0.4533	0.87527954		
+	0.4534	0.89798489		
+	0.4535	0.89234712		
+	0.4536	0.89474958		
+	0.4537	0.89718319		
+	0.4538	0.90433579		
+	0.4539	0.90261376		
+	0.454	0.88703673		
+	0.4541	0.88949036		
+	0.4542	0.88366462		
+	0.4543	0.88831168		
+	0.4544	0.88830944		
+	0.4545	0.88785643		
+	0.4546	0.87370833		
+	0.4547	0.86886571		
+	0.4548	0.86085213		
+	0.4549	0.85927616		
+	0.455	0.85130622		
+	0.4551	0.84818822		
+	0.4552	0.8575061		
+	0.4553	0.8609639		
+	0.4554	0.84654875		
+	0.4555	0.84756912		
+	0.4556	0.84644485		
+	0.4557	0.84650534		
+	0.4558	0.84262852		
+	0.4559	0.85629206		
+	0.456	0.85906293		
+	0.4561	0.87112625		
+	0.4562	0.88453088		
+	0.4563	0.88857012		
+	0.4564	0.89550374		
+	0.4565	0.89731583		
+	0.4566	0.89154807		
+	0.4567	0.88839179		
+	0.4568	0.90427117		
+	0.4569	0.8961241		
+	0.457	0.89048523		
+	0.4571	0.90225027		
+	0.4572	0.90658204		
+	0.4573	0.89816497		
+	0.4574	0.8891171		
+	0.4575	0.89002674		
+	0.4576	0.90097163		
+	0.4577	0.90660047		
+	0.4578	0.90000824		
+	0.4579	0.89581149		
+	0.458	0.89994768		
+	0.4581	0.91113062		
+	0.4582	0.89928456		
+	0.4583	0.91743803		
+	0.4584	0.91387728		
+	0.4585	0.91065302		
+	0.4586	0.92784255		
+	0.4587	0.93561681		
+	0.4588	0.93060809		
+	0.4589	0.94235809		
+	0.459	0.95177588		
+	0.4591	0.9703066		
+	0.4592	0.9872621		
+	0.4593	0.99154054		
+	0.4594	1.0002438		
+	0.4595	0.9880753		
+	0.4596	0.99258583		
+	0.4597	0.99462359		
+	0.4598	0.99730545		
+	0.4599	0.99924587		
+	0.46	0.99504807		
+	0.4601	0.99915642		
+	0.4602	0.99339891		
+	0.4603	0.98238064		
+	0.4604	0.98812914		
+	0.4605	0.98780649		
+	0.4606	0.96626563		
+	0.4607	0.9729007		
+	0.4608	0.96886814		
+	0.4609	0.97502731		
+	0.461	0.96849133		
+	0.4611	0.96318718		
+	0.4612	0.95953512		
+	0.4613	0.95455522		
+	0.4614	0.94741653		
+	0.4615	0.95527069		
+	0.4616	0.9488998		
+	0.4617	0.96488264		
+	0.4618	0.96740266		
+	0.4619	0.97416851		
+	0.462	0.98960478		
+	0.4621	0.98485766		
+	0.4622	1.0026745		
+	0.4623	1.0123887		
+	0.4624	1.0154537		
+	0.4625	1.0167131		
+	0.4626	1.012469		
+	0.4627	0.99453097		
+	0.4628	0.99652333		
+	0.4629	0.99207237		
+	0.463	1.0070399		
+	0.4631	1.0042184		
+	0.4632	0.99678638		
+	0.4633	0.97813848		
+	0.4634	0.97376976		
+	0.4635	0.97751841		
+	0.4636	0.98134524		
+	0.4637	0.97496		
+	0.4638	0.95819742		
+	0.4639	0.9511201		
+	0.464	0.95946109		
+	0.4641	0.93948753		
+	0.4642	0.94535545		
+	0.4643	0.92350386		
+	0.4644	0.91908136		
+	0.4645	0.91281912		
+	0.4646	0.90102505		
+	0.4647	0.90511007		
+	0.4648	0.91695666		
+	0.4649	0.91195536		
+	0.465	0.91352676		
+	0.4651	0.92914739		
+	0.4652	0.93454576		
+	0.4653	0.91855629		
+	0.4654	0.91610788		
+	0.4655	0.92147134		
+	0.4656	0.91698984		
+	0.4657	0.91068573		
+	0.4658	0.90592753		
+	0.4659	0.89698947		
+	0.466	0.89834863		
+	0.4661	0.87989104		
+	0.4662	0.87120847		
+	0.4663	0.87309563		
+	0.4664	0.86502723		
+	0.4665	0.86501878		
+	0.4666	0.86735363		
+	0.4667	0.8569413		
+	0.4668	0.85135186		
+	0.4669	0.85284635		
+	0.467	0.8438999		
+	0.4671	0.83804015		
+	0.4672	0.84238852		
+	0.4673	0.84816466		
+	0.4674	0.83200489		
+	0.4675	0.83615083		
+	0.4676	0.83629253		
+	0.4677	0.84856551		
+	0.4678	0.85809051		
+	0.4679	0.87826686		
+	0.468	0.88834969		
+	0.4681	0.87673029		
+	0.4682	0.89473785		
+	0.4683	0.88780268		
+	0.4684	0.88970915		
+	0.4685	0.88697971		
+	0.4686	0.88139563		
+	0.4687	0.88002038		
+	0.4688	0.87767127		
+	0.4689	0.88648216		
+	0.469	0.8834193		
+	0.4691	0.86846051		
+	0.4692	0.87577903		
+	0.4693	0.8675099		
+	0.4694	0.86782878		
+	0.4695	0.85455409		
+	0.4696	0.84559783		
+	0.4697	0.85391695		
+	0.4698	0.83668228		
+	0.4699	0.83856811		
+	0.47	0.8386608		
+	0.4701	0.84544507		
+	0.4702	0.84393927		
+	0.4703	0.84690951		
+	0.4704	0.84360732		
+	0.4705	0.83315197		
+	0.4706	0.84679853		
+	0.4707	0.85852055		
+	0.4708	0.87081014		
+	0.4709	0.88113516		
+	0.471	0.88260917		
+	0.4711	0.89095798		
+	0.4712	0.8914848		
+	0.4713	0.8809341		
+	0.4714	0.88975549		
+	0.4715	0.87702489		
+	0.4716	0.88452273		
+	0.4717	0.8877062		
+	0.4718	0.87494013		
+	0.4719	0.86802758		
+	0.472	0.87322419		
+	0.4721	0.85891718		
+	0.4722	0.85864238		
+	0.4723	0.86475474		
+	0.4724	0.85255583		
+	0.4725	0.85988772		
+	0.4726	0.84165088		
+	0.4727	0.85316984		
+	0.4728	0.84817372		
+	0.4729	0.84172134		
+	0.473	0.84066781		
+	0.4731	0.84375504		
+	0.4732	0.84744157		
+	0.4733	0.84495837		
+	0.4734	0.84159393		
+	0.4735	0.84751536		
+	0.4736	0.86504469		
+	0.4737	0.8772164		
+	0.4738	0.8960199		
+	0.4739	0.90480299		
+	0.474	0.90475557		
+	0.4741	0.91682599		
+	0.4742	0.91371212		
+	0.4743	0.92489976		
+	0.4744	0.92777201		
+	0.4745	0.9412609		
+	0.4746	0.93595751		
+	0.4747	0.94441849		
+	0.4748	0.94353568		
+	0.4749	0.95628041		
+	0.475	0.94285372		
+	0.4751	0.95713096		
+	0.4752	0.95143042		
+	0.4753	0.96082623		
+	0.4754	0.94273321		
+	0.4755	0.95679225		
+	0.4756	0.94778064		
+	0.4757	0.94069416		
+	0.4758	0.9515923		
+	0.4759	0.95013308		
+	0.476	0.93691893		
+	0.4761	0.93859381		
+	0.4762	0.93672504		
+	0.4763	0.93552233		
+	0.4764	0.94883093		
+	0.4765	0.94756866		
+	0.4766	0.95923259		
+	0.4767	0.97194358		
+	0.4768	0.98447119		
+	0.4769	0.98731812		
+	0.477	1.0034247		
+	0.4771	1.0052368		
+	0.4772	0.98737046		
+	0.4773	1.0007379		
+	0.4774	0.98899458		
+	0.4775	0.98671487		
+	0.4776	0.99146735		
+	0.4777	0.99250673		
+	0.4778	0.99183467		
+	0.4779	0.98120598		
+	0.478	0.97065242		
+	0.4781	0.98037109		
+	0.4782	0.96861005		
+	0.4783	0.97249804		
+	0.4784	0.96020052		
+	0.4785	0.96056888		
+	0.4786	0.96009486		
+	0.4787	0.95382312		
+	0.4788	0.95099811		
+	0.4789	0.9471651		
+	0.479	0.93771278		
+	0.4791	0.94437103		
+	0.4792	0.93801077		
+	0.4793	0.94691831		
+	0.4794	0.95334091		
+	0.4795	0.97749431		
+	0.4796	0.97576145		
+	0.4797	0.99024767		
+	0.4798	0.99209219		
+	0.4799	0.98895071		
+	0.48	1.0030714		
+	0.4801	0.98144053		
+	0.4802	0.97802689		
+	0.4803	0.98221381		
+	0.4804	0.97436406		
+	0.4805	0.95227884		
+	0.4806	0.95584818		
+	0.4807	0.93881687		
+	0.4808	0.92277255		
+	0.4809	0.92297154		
+	0.481	0.91330982		
+	0.4811	0.90010466		
+	0.4812	0.894614		
+	0.4813	0.87570531		
+	0.4814	0.86356923		
+	0.4815	0.86831667		
+	0.4816	0.8665309		
+	0.4817	0.85335022		
+	0.4818	0.84069876		
+	0.4819	0.84941209		
+	0.482	0.83578307		
+	0.4821	0.84287875		
+	0.4822	0.83203622		
+	0.4823	0.8510304		
+	0.4824	0.85311127		
+	0.4825	0.85378926		
+	0.4826	0.87547132		
+	0.4827	0.87223765		
+	0.4828	0.88490161		
+	0.4829	0.88238571		
+	0.483	0.88027417		
+	0.4831	0.88522549		
+	0.4832	0.8712672		
+	0.4833	0.87328567		
+	0.4834	0.87411477		
+	0.4835	0.87696741		
+	0.4836	0.85551431		
+	0.4837	0.85666058		
+	0.4838	0.85239374		
+	0.4839	0.84490735		
+	0.484	0.85130527		
+	0.4841	0.85316371		
+	0.4842	0.84740852		
+	0.4843	0.84008128		
+	0.4844	0.84097239		
+	0.4845	0.83680564		
+	0.4846	0.83508855		
+	0.4847	0.83973274		
+	0.4848	0.83025193		
+	0.4849	0.81829308		
+	0.485	0.82263436		
+	0.4851	0.83624835		
+	0.4852	0.83860246		
+	0.4853	0.84013078		
+	0.4854	0.84970186		
+	0.4855	0.86604151		
+	0.4856	0.8701595		
+	0.4857	0.87120404		
+	0.4858	0.8801303		
+	0.4859	0.87507811		
+	0.486	0.88577273		
+	0.4861	0.86706839		
+	0.4862	0.88262282		
+	0.4863	0.8753919		
+	0.4864	0.86335849		
+	0.4865	0.8661769		
+	0.4866	0.8649873		
+	0.4867	0.86273088		
+	0.4868	0.85635367		
+	0.4869	0.84466623		
+	0.487	0.84728357		
+	0.4871	0.83961645		
+	0.4872	0.84133477		
+	0.4873	0.84275685		
+	0.4874	0.83719916		
+	0.4875	0.83059323		
+	0.4876	0.83439036		
+	0.4877	0.83130365		
+	0.4878	0.83188798		
+	0.4879	0.82052796		
+	0.488	0.8370768		
+	0.4881	0.84262151		
+	0.4882	0.83846199		
+	0.4883	0.85312286		
+	0.4884	0.86034922		
+	0.4885	0.86341073		
+	0.4886	0.86766109		
+	0.4887	0.88630528		
+	0.4888	0.87181715		
+	0.4889	0.87884669		
+	0.489	0.87488046		
+	0.4891	0.87637573		
+	0.4892	0.87703002		
+	0.4893	0.87810029		
+	0.4894	0.8703392		
+	0.4895	0.85576672		
+	0.4896	0.86699215		
+	0.4897	0.86356522		
+	0.4898	0.86103189		
+	0.4899	0.84957043		
+	0.49	0.85562602		
+	0.4901	0.8519825		
+	0.4902	0.8529811		
+	0.4903	0.85421946		
+	0.4904	0.85623906		
+	0.4905	0.86880625		
+	0.4906	0.86608979		
+	0.4907	0.87183132		
+	0.4908	0.89250571		
+	0.4909	0.89700403		
+	0.491	0.89464278		
+	0.4911	0.92112072		
+	0.4912	0.94189109		
+	0.4913	0.94592807		
+	0.4914	0.95262731		
+	0.4915	0.96630244		
+	0.4916	0.96838953		
+	0.4917	0.98493881		
+	0.4918	0.98487476		
+	0.4919	0.96729693		
+	0.492	0.97750637		
+	0.4921	0.96946368		
+	0.4922	0.97148255		
+	0.4923	0.9771554		
+	0.4924	0.97120098		
+	0.4925	0.97177204		
+	0.4926	0.96610927		
+	0.4927	0.94696988		
+	0.4928	0.95490741		
+	0.4929	0.94728949		
+	0.493	0.95580764		
+	0.4931	0.93540356		
+	0.4932	0.94262656		
+	0.4933	0.94100788		
+	0.4934	0.9462717		
+	0.4935	0.93008634		
+	0.4936	0.93072912		
+	0.4937	0.94394366		
+	0.4938	0.94500193		
+	0.4939	0.94798418		
+	0.494	0.95137586		
+	0.4941	0.94911485		
+	0.4942	0.96357872		
+	0.4943	0.97150627		
+	0.4944	0.98847897		
+	0.4945	0.98783775		
+	0.4946	0.99367533		
+	0.4947	0.9887591		
+	0.4948	0.98762278		
+	0.4949	0.98166423		
+	0.495	0.97388844		
+	0.4951	0.97719309		
+	0.4952	0.98433063		
+	0.4953	0.96752624		
+	0.4954	0.97015831		
+	0.4955	0.97356307		
+	0.4956	0.96813206		
+	0.4957	0.95232802		
+	0.4958	0.95973627		
+	0.4959	0.9544306		
+	0.496	0.95427038		
+	0.4961	0.94628998		
+	0.4962	0.93779031		
+	0.4963	0.92298961		
+	0.4964	0.92786571		
+	0.4965	0.92936953		
+	0.4966	0.91815194		
+	0.4967	0.90867024		
+	0.4968	0.89087641		
+	0.4969	0.8941514		
+	0.497	0.9029773		
+	0.4971	0.89845812		
+	0.4972	0.9033173		
+	0.4973	0.90289958		
+	0.4974	0.90337168		
+	0.4975	0.91657163		
+	0.4976	0.90060446		
+	0.4977	0.88807022		
+	0.4978	0.89872445		
+	0.4979	0.8913238		
+	0.498	0.88884377		
+	0.4981	0.86857919		
+	0.4982	0.86836503		
+	0.4983	0.85506743		
+	0.4984	0.85465452		
+	0.4985	0.8486016		
+	0.4986	0.83908394		
+	0.4987	0.84165474		
+	0.4988	0.82628775		
+	0.4989	0.82946372		
+	0.499	0.8278463		
+	0.4991	0.83295571		
+	0.4992	0.82539018		
+	0.4993	0.8196183		
+	0.4994	0.82442526		
+	0.4995	0.82173625		
+	0.4996	0.81458595		
+	0.4997	0.81613753		
+	0.4998	0.82721637		
+	0.4999	0.82662189		
+	0.5	0.83608077		
+	0.5001	0.86010015		
+	0.5002	0.85362067		
+	0.5003	0.86212958		
+	0.5004	0.87212788		
+	0.5005	0.87210475		
+	0.5006	0.86722762		
+	0.5007	0.86003132		
+	0.5008	0.86703951		
+	0.5009	0.85501605		
+	0.501	0.85468534		
+	0.5011	0.8630337		
+	0.5012	0.85511719		
+	0.5013	0.85799439		
+	0.5014	0.84493508		
+	0.5015	0.83461701		
+	0.5016	0.83524049		
+	0.5017	0.84065751		
+	0.5018	0.82734897		
+	0.5019	0.81940039		
+	0.502	0.82665942		
+	0.5021	0.82188755		
+	0.5022	0.8256144		
+	0.5023	0.82643434		
+	0.5024	0.80826996		
+	0.5025	0.81634478		
+	0.5026	0.82251859		
+	0.5027	0.8267175		
+	0.5028	0.83764882		
+	0.5029	0.844819		
+	0.503	0.84452777		
+	0.5031	0.86156053		
+	0.5032	0.86879336		
+	0.5033	0.86726995		
+	0.5034	0.86904133		
+	0.5035	0.87510801		
+	0.5036	0.85702231		
+	0.5037	0.86283655		
+	0.5038	0.86457818		
+	0.5039	0.85409986		
+	0.504	0.85363199		
+	0.5041	0.85628709		
+	0.5042	0.84956313		
+	0.5043	0.84521932		
+	0.5044	0.8479687		
+	0.5045	0.84097257		
+	0.5046	0.82718308		
+	0.5047	0.83776814		
+	0.5048	0.82676205		
+	0.5049	0.81848002		
+	0.505	0.82853833		
+	0.5051	0.82709457		
+	0.5052	0.80763603		
+	0.5053	0.81070622		
+	0.5054	0.81550296		
+	0.5055	0.80727542		
+	0.5056	0.82407358		
+	0.5057	0.81857517		
+	0.5058	0.83445949		
+	0.5059	0.85210616		
+	0.506	0.86846235		
+	0.5061	0.86533386		
+	0.5062	0.88183646		
+	0.5063	0.89291796		
+	0.5064	0.89312819		
+	0.5065	0.89502607		
+	0.5066	0.89782089		
+	0.5067	0.90286211		
+	0.5068	0.90916193		
+	0.5069	0.90468054		
+	0.507	0.91147265		
+	0.5071	0.90918857		
+	0.5072	0.90795635		
+	0.5073	0.92321742		
+	0.5074	0.91997694		
+	0.5075	0.91167395		
+	0.5076	0.92506751		
+	0.5077	0.91593041		
+	0.5078	0.92594806		
+	0.5079	0.92931158		
+	0.508	0.91930359		
+	0.5081	0.91679051		
+	0.5082	0.90943534		
+	0.5083	0.90881167		
+	0.5084	0.9192177		
+	0.5085	0.91859158		
+	0.5086	0.93382277		
+	0.5087	0.93827355		
+	0.5088	0.95490384		
+	0.5089	0.95558344		
+	0.509	0.97179869		
+	0.5091	0.97360447		
+	0.5092	0.96623079		
+	0.5093	0.97361942		
+	0.5094	0.96737054		
+	0.5095	0.97415204		
+	0.5096	0.95940747		
+	0.5097	0.9703849		
+	0.5098	0.97049747		
+	0.5099	0.95843696		
+	0.51	0.95681542		
+	0.5101	0.94555189		
+	0.5102	0.95252114		
+	0.5103	0.93981931		
+	0.5104	0.94266217		
+	0.5105	0.93928033		
+	0.5106	0.93953305		
+	0.5107	0.92374776		
+	0.5108	0.93415497		
+	0.5109	0.93377977		
+	0.511	0.93037772		
+	0.5111	0.93355523		
+	0.5112	0.93112229		
+	0.5113	0.92560049		
+	0.5114	0.92743768		
+	0.5115	0.92483416		
+	0.5116	0.93870003		
+	0.5117	0.9505788		
+	0.5118	0.95667822		
+	0.5119	0.97263752		
+	0.512	0.97874075		
+	0.5121	0.98051612		
+	0.5122	0.97680024		
+	0.5123	0.97445321		
+	0.5124	0.97119394		
+	0.5125	0.96287853		
+	0.5126	0.96028814		
+	0.5127	0.96081807		
+	0.5128	0.95028323		
+	0.5129	0.93913455		
+	0.513	0.91343935		
+	0.5131	0.91333391		
+	0.5132	0.88779287		
+	0.5133	0.87845612		
+	0.5134	0.88490037		
+	0.5135	0.86490254		
+	0.5136	0.86602553		
+	0.5137	0.84796677		
+	0.5138	0.8527482		
+	0.5139	0.83083102		
+	0.514	0.84394526		
+	0.5141	0.82884212		
+	0.5142	0.83570795		
+	0.5143	0.83347413		
+	0.5144	0.82920301		
+	0.5145	0.83075162		
+	0.5146	0.84246294		
+	0.5147	0.85142698		
+	0.5148	0.85954284		
+	0.5149	0.85912957		
+	0.515	0.85550343		
+	0.5151	0.86758741		
+	0.5152	0.85446402		
+	0.5153	0.84997523		
+	0.5154	0.85150794		
+	0.5155	0.85101044		
+	0.5156	0.85785549		
+	0.5157	0.85278533		
+	0.5158	0.8506045		
+	0.5159	0.84042499		
+	0.516	0.82774019		
+	0.5161	0.82512373		
+	0.5162	0.82186147		
+	0.5163	0.83110906		
+	0.5164	0.82086091		
+	0.5165	0.82365511		
+	0.5166	0.81158351		
+	0.5167	0.80829231		
+	0.5168	0.81350905		
+	0.5169	0.81283308		
+	0.517	0.80377234		
+	0.5171	0.81088571		
+	0.5172	0.79894847		
+	0.5173	0.80674017		
+	0.5174	0.82013357		
+	0.5175	0.82621989		
+	0.5176	0.83397865		
+	0.5177	0.85597022		
+	0.5178	0.84907774		
+	0.5179	0.84701521		
+	0.518	0.86432867		
+	0.5181	0.85700562		
+	0.5182	0.85431752		
+	0.5183	0.85416317		
+	0.5184	0.85696799		
+	0.5185	0.85061215		
+	0.5186	0.8397101		
+	0.5187	0.83502897		
+	0.5188	0.84745258		
+	0.5189	0.83845561		
+	0.519	0.8244287		
+	0.5191	0.8215826		
+	0.5192	0.8176869		
+	0.5193	0.81042367		
+	0.5194	0.81477219		
+	0.5195	0.81920674		
+	0.5196	0.82052221		
+	0.5197	0.80701547		
+	0.5198	0.81583796		
+	0.5199	0.80139171		
+	0.52	0.79540709		
+	0.5201	0.80692941		
+	0.5202	0.8054152		
+	0.5203	0.8072685		
+	0.5204	0.81655742		
+	0.5205	0.83452978		
+	0.5206	0.85232301		
+	0.5207	0.84250091		
+	0.5208	0.86491416		
+	0.5209	0.86309359		
+	0.521	0.85481084		
+	0.5211	0.85098577		
+	0.5212	0.85232108		
+	0.5213	0.84807372		
+	0.5214	0.85255372		
+	0.5215	0.853502		
+	0.5216	0.83962227		
+	0.5217	0.83477906		
+	0.5218	0.83167901		
+	0.5219	0.82841903		
+	0.522	0.82308417		
+	0.5221	0.83020917		
+	0.5222	0.81813349		
+	0.5223	0.8214909		
+	0.5224	0.83740096		
+	0.5225	0.8323764		
+	0.5226	0.84151609		
+	0.5227	0.826372		
+	0.5228	0.83728108		
+	0.5229	0.85154794		
+	0.523	0.84340348		
+	0.5231	0.84740417		
+	0.5232	0.85797083		
+	0.5233	0.87515855		
+	0.5234	0.90725924		
+	0.5235	0.91593553		
+	0.5236	0.92379195		
+	0.5237	0.94205157		
+	0.5238	0.94944257		
+	0.5239	0.94941777		
+	0.524	0.95613177		
+	0.5241	0.94311675		
+	0.5242	0.95160908		
+	0.5243	0.94316049		
+	0.5244	0.95237294		
+	0.5245	0.95011174		
+	0.5246	0.9365024		
+	0.5247	0.94310653		
+	0.5248	0.92555362		
+	0.5249	0.927294		
+	0.525	0.92715947		
+	0.5251	0.93104128		
+	0.5252	0.91248201		
+	0.5253	0.92892335		
+	0.5254	0.91950787		
+	0.5255	0.90691584		
+	0.5256	0.91451364		
+	0.5257	0.90590968		
+	0.5258	0.90910065		
+	0.5259	0.90831466		
+	0.526	0.91903888		
+	0.5261	0.9109399		
+	0.5262	0.91835929		
+	0.5263	0.94138778		
+	0.5264	0.9404035		
+	0.5265	0.95649827		
+	0.5266	0.95426722		
+	0.5267	0.97016055		
+	0.5268	0.97183033		
+	0.5269	0.96156338		
+	0.527	0.9558197		
+	0.5271	0.95026401		
+	0.5272	0.94991769		
+	0.5273	0.95744567		
+	0.5274	0.96004537		
+	0.5275	0.95522879		
+	0.5276	0.94905101		
+	0.5277	0.94684988		
+	0.5278	0.94773017		
+	0.5279	0.93888456		
+	0.528	0.93028941		
+	0.5281	0.93267883		
+	0.5282	0.92483812		
+	0.5283	0.92457954		
+	0.5284	0.92209197		
+	0.5285	0.92407294		
+	0.5286	0.90149186		
+	0.5287	0.91140435		
+	0.5288	0.90789005		
+	0.5289	0.89194863		
+	0.529	0.88982567		
+	0.5291	0.88772626		
+	0.5292	0.88848756		
+	0.5293	0.90674809		
+	0.5294	0.89943293		
+	0.5295	0.9075374		
+	0.5296	0.90825887		
+	0.5297	0.89167238		
+	0.5298	0.89542931		
+	0.5299	0.8786159		
+	0.53	0.87625394		
+	0.5301	0.86976913		
+	0.5302	0.87526809		
+	0.5303	0.85127604		
+	0.5304	0.85310813		
+	0.5305	0.84757628		
+	0.5306	0.84008623		
+	0.5307	0.84312417		
+	0.5308	0.81956953		
+	0.5309	0.81975737		
+	0.531	0.8221009		
+	0.5311	0.81346454		
+	0.5312	0.80440714		
+	0.5313	0.80355774		
+	0.5314	0.79746026		
+	0.5315	0.80353771		
+	0.5316	0.79741075		
+	0.5317	0.79702117		
+	0.5318	0.80232621		
+	0.5319	0.80601541		
+	0.532	0.81459886		
+	0.5321	0.80901081		
+	0.5322	0.8228812		
+	0.5323	0.83240216		
+	0.5324	0.84154262		
+	0.5325	0.84765485		
+	0.5326	0.85111112		
+	0.5327	0.84462602		
+	0.5328	0.84891806		
+	0.5329	0.83731583		
+	0.533	0.83736655		
+	0.5331	0.84560474		
+	0.5332	0.84486442		
+	0.5333	0.83761164		
+	0.5334	0.82146446		
+	0.5335	0.83172839		
+	0.5336	0.82837599		
+	0.5337	0.81901687		
+	0.5338	0.8153098		
+	0.5339	0.8181395		
+	0.534	0.81573771		
+	0.5341	0.81277107		
+	0.5342	0.80352019		
+	0.5343	0.79091115		
+	0.5344	0.80231303		
+	0.5345	0.79585671		
+	0.5346	0.79679262		
+	0.5347	0.79044233		
+	0.5348	0.7968645		
+	0.5349	0.79874899		
+	0.535	0.8050985		
+	0.5351	0.82833127		
+	0.5352	0.82498753		
+	0.5353	0.84226793		
+	0.5354	0.83824343		
+	0.5355	0.85682566		
+	0.5356	0.84759051		
+	0.5357	0.84803854		
+	0.5358	0.84558994		
+	0.5359	0.83734087		
+	0.536	0.84135821		
+	0.5361	0.8357939		
+	0.5362	0.84147224		
+	0.5363	0.83937985		
+	0.5364	0.83252402		
+	0.5365	0.81507282		
+	0.5366	0.81706025		
+	0.5367	0.8244515		
+	0.5368	0.81884346		
+	0.5369	0.80027007		
+	0.537	0.7975423		
+	0.5371	0.80792831		
+	0.5372	0.79370866		
+	0.5373	0.79759029		
+	0.5374	0.7919937		
+	0.5375	0.79173363		
+	0.5376	0.78559293		
+	0.5377	0.7979876		
+	0.5378	0.7942447		
+	0.5379	0.80426812		
+	0.538	0.82902563		
+	0.5381	0.8286015		
+	0.5382	0.83362208		
+	0.5383	0.84116407		
+	0.5384	0.85486528		
+	0.5385	0.86358757		
+	0.5386	0.85609331		
+	0.5387	0.86200253		
+	0.5388	0.86971181		
+	0.5389	0.86529358		
+	0.539	0.86503168		
+	0.5391	0.87885589		
+	0.5392	0.86564913		
+	0.5393	0.88203978		
+	0.5394	0.87769115		
+	0.5395	0.88429619		
+	0.5396	0.87485477		
+	0.5397	0.89412787		
+	0.5398	0.88321909		
+	0.5399	0.88246791		
+	0.54	0.89456665		
+	0.5401	0.89998857		
+	0.5402	0.89233215		
+	0.5403	0.90220309		
+	0.5404	0.88461668		
+	0.5405	0.9022345		
+	0.5406	0.88853753		
+	0.5407	0.89859133		
+	0.5408	0.90615457		
+	0.5409	0.92360713		
+	0.541	0.93566376		
+	0.5411	0.94098256		
+	0.5412	0.94977049		
+	0.5413	0.95634791		
+	0.5414	0.955487		
+	0.5415	0.94501972		
+	0.5416	0.95978483		
+	0.5417	0.95044492		
+	0.5418	0.95577711		
+	0.5419	0.94095087		
+	0.542	0.95245417		
+	0.5421	0.94835222		
+	0.5422	0.94619586		
+	0.5423	0.94333493		
+	0.5424	0.93800487		
+	0.5425	0.92025881		
+	0.5426	0.9125595		
+	0.5427	0.92783203		
+	0.5428	0.91358718		
+	0.5429	0.90211126		
+	0.543	0.90252052		
+	0.5431	0.90857525		
+	0.5432	0.90860672		
+	0.5433	0.90482977		
+	0.5434	0.89361908		
+	0.5435	0.89703069		
+	0.5436	0.91589445		
+	0.5437	0.91547901		
+	0.5438	0.92847214		
+	0.5439	0.94358181		
+	0.544	0.94669868		
+	0.5441	0.94864003		
+	0.5442	0.9467865		
+	0.5443	0.96122103		
+	0.5444	0.95072019		
+	0.5445	0.96038842		
+	0.5446	0.94796066		
+	0.5447	0.95166306		
+	0.5448	0.95165709		
+	0.5449	0.93852159		
+	0.545	0.92488783		
+	0.5451	0.93357026		
+	0.5452	0.92558672		
+	0.5453	0.90831574		
+	0.5454	0.88296741		
+	0.5455	0.88878708		
+	0.5456	0.86102969		
+	0.5457	0.86118034		
+	0.5458	0.85081801		
+	0.5459	0.83855333		
+	0.546	0.8341364		
+	0.5461	0.830894		
+	0.5462	0.82425897		
+	0.5463	0.81946503		
+	0.5464	0.82186649		
+	0.5465	0.81711876		
+	0.5466	0.82278691		
+	0.5467	0.81893524		
+	0.5468	0.83957722		
+	0.5469	0.84271433		
+	0.547	0.83875786		
+	0.5471	0.84977002		
+	0.5472	0.85232184		
+	0.5473	0.83719798		
+	0.5474	0.85064265		
+	0.5475	0.84524801		
+	0.5476	0.84432547		
+	0.5477	0.83974587		
+	0.5478	0.8391485		
+	0.5479	0.81939496		
+	0.548	0.82698324		
+	0.5481	0.82401449		
+	0.5482	0.81953861		
+	0.5483	0.81190563		
+	0.5484	0.80163169		
+	0.5485	0.80245526		
+	0.5486	0.79221831		
+	0.5487	0.80034361		
+	0.5488	0.79382665		
+	0.5489	0.79070928		
+	0.549	0.79640123		
+	0.5491	0.79555557		
+	0.5492	0.7916179		
+	0.5493	0.77828362		
+	0.5494	0.79089739		
+	0.5495	0.78421486		
+	0.5496	0.79864368		
+	0.5497	0.81711816		
+	0.5498	0.82117199		
+	0.5499	0.83583205		
+	0.55	0.84181655		
+	0.5501	0.84760993		
+	0.5502	0.83029144		
+	0.5503	0.833825		
+	0.5504	0.83063		
+	0.5505	0.84242066		
+	0.5506	0.8310206		
+	0.5507	0.83256729		
+	0.5508	0.82461027		
+	0.5509	0.82685607		
+	0.551	0.82877113		
+	0.5511	0.81900647		
+	0.5512	0.81940306		
+	0.5513	0.8044752		
+	0.5514	0.80677244		
+	0.5515	0.79683167		
+	0.5516	0.79934023		
+	0.5517	0.80406327		
+	0.5518	0.78503653		
+	0.5519	0.79777622		
+	0.552	0.79915011		
+	0.5521	0.79325851		
+	0.5522	0.78440433		
+	0.5523	0.79045502		
+	0.5524	0.79613325		
+	0.5525	0.80157406		
+	0.5526	0.80608326		
+	0.5527	0.8299614		
+	0.5528	0.83711773		
+	0.5529	0.83689216		
+	0.553	0.8354092		
+	0.5531	0.83671824		
+	0.5532	0.83181311		
+	0.5533	0.83569843		
+	0.5534	0.8368752		
+	0.5535	0.83984916		
+	0.5536	0.82416772		
+	0.5537	0.83516396		
+	0.5538	0.82664441		
+	0.5539	0.82672573		
+	0.554	0.8247117		
+	0.5541	0.81112459		
+	0.5542	0.80024423		
+	0.5543	0.80429942		
+	0.5544	0.79919935		
+	0.5545	0.81019294		
+	0.5546	0.80041499		
+	0.5547	0.80364933		
+	0.5548	0.80949636		
+	0.5549	0.81145213		
+	0.555	0.8170087		
+	0.5551	0.81450852		
+	0.5552	0.81142679		
+	0.5553	0.83750465		
+	0.5554	0.84810327		
+	0.5555	0.86225826		
+	0.5556	0.87959327		
+	0.5557	0.878664		
+	0.5558	0.91009885		
+	0.5559	0.91831163		
+	0.556	0.91508427		
+	0.5561	0.92444263		
+	0.5562	0.92430223		
+	0.5563	0.92046272		
+	0.5564	0.93491067		
+	0.5565	0.93566979		
+	0.5566	0.93758014		
+	0.5567	0.92644242		
+	0.5568	0.92598745		
+	0.5569	0.91740097		
+	0.557	0.9165762		
+	0.5571	0.91149596		
+	0.5572	0.90991471		
+	0.5573	0.89660108		
+	0.5574	0.91006974		
+	0.5575	0.91008913		
+	0.5576	0.90302609		
+	0.5577	0.90214005		
+	0.5578	0.89422109		
+	0.5579	0.89378823		
+	0.558	0.88711082		
+	0.5581	0.88960138		
+	0.5582	0.89296254		
+	0.5583	0.89575399		
+	0.5584	0.91319059		
+	0.5585	0.93251797		
+	0.5586	0.93358674		
+	0.5587	0.93680507		
+	0.5588	0.94668346		
+	0.5589	0.95810461		
+	0.559	0.95719922		
+	0.5591	0.94756261		
+	0.5592	0.93901805		
+	0.5593	0.9392834		
+	0.5594	0.94798151		
+	0.5595	0.92990922		
+	0.5596	0.92945389		
+	0.5597	0.93042784		
+	0.5598	0.92829163		
+	0.5599	0.92788554		
+	0.56	0.91998733		
+	0.5601	0.91032775		
+	0.5602	0.91647454		
+	0.5603	0.915402		
+	0.5604	0.9118142		
+	0.5605	0.91158329		
+	0.5606	0.9088341		
+	0.5607	0.91016673		
+	0.5608	0.8959057		
+	0.5609	0.88683738		
+	0.561	0.89188175		
+	0.5611	0.89073915		
+	0.5612	0.89464561		
+	0.5613	0.91075562		
+	0.5614	0.9054076		
+	0.5615	0.91795198		
+	0.5616	0.91287125		
+	0.5617	0.9148566		
+	0.5618	0.89813031		
+	0.5619	0.89024788		
+	0.562	0.88345346		
+	0.5621	0.89055787		
+	0.5622	0.88327363		
+	0.5623	0.86518332		
+	0.5624	0.8638693		
+	0.5625	0.85755718		
+	0.5626	0.84841443		
+	0.5627	0.84447089		
+	0.5628	0.83832311		
+	0.5629	0.83359049		
+	0.563	0.82719037		
+	0.5631	0.80220779		
+	0.5632	0.81417526		
+	0.5633	0.80080382		
+	0.5634	0.80178425		
+	0.5635	0.79537149		
+	0.5636	0.7850454		
+	0.5637	0.7924424		
+	0.5638	0.79085284		
+	0.5639	0.78947178		
+	0.564	0.78009946		
+	0.5641	0.78166787		
+	0.5642	0.79810412		
+	0.5643	0.80954491		
+	0.5644	0.810529		
+	0.5645	0.82587318		
+	0.5646	0.83449839		
+	0.5647	0.84173183		
+	0.5648	0.83192261		
+	0.5649	0.83270641		
+	0.565	0.82658292		
+	0.5651	0.82927756		
+	0.5652	0.83539448		
+	0.5653	0.81915462		
+	0.5654	0.82511849		
+	0.5655	0.81953294		
+	0.5656	0.81030397		
+	0.5657	0.81549547		
+	0.5658	0.79977073		
+	0.5659	0.79659991		
+	0.566	0.79232058		
+	0.5661	0.80253923		
+	0.5662	0.79375615		
+	0.5663	0.78413371		
+	0.5664	0.78450156		
+	0.5665	0.78395409		
+	0.5666	0.79209981		
+	0.5667	0.78428535		
+	0.5668	0.78179762		
+	0.5669	0.77751493		
+	0.567	0.77889462		
+	0.5671	0.78572101		
+	0.5672	0.79997679		
+	0.5673	0.82046262		
+	0.5674	0.81679051		
+	0.5675	0.83039412		
+	0.5676	0.83488159		
+	0.5677	0.84340235		
+	0.5678	0.84274193		
+	0.5679	0.82817906		
+	0.568	0.82769439		
+	0.5681	0.82258722		
+	0.5682	0.82709456		
+	0.5683	0.8331487		
+	0.5684	0.82219339		
+	0.5685	0.80669871		
+	0.5686	0.82067588		
+	0.5687	0.80845714		
+	0.5688	0.80381162		
+	0.5689	0.80626556		
+	0.569	0.80521498		
+	0.5691	0.80184472		
+	0.5692	0.78897056		
+	0.5693	0.79588536		
+	0.5694	0.78439826		
+	0.5695	0.78411392		
+	0.5696	0.78148701		
+	0.5697	0.78388148		
+	0.5698	0.7906521		
+	0.5699	0.77956794		
+	0.57	0.78822466		
+	0.5701	0.80831769		
+	0.5702	0.81497335		
+	0.5703	0.82580502		
+	0.5704	0.82790231		
+	0.5705	0.83351221		
+	0.5706	0.83987665		
+	0.5707	0.83017096		
+	0.5708	0.83103866		
+	0.5709	0.84027304		
+	0.571	0.83356966		
+	0.5711	0.83443112		
+	0.5712	0.85103225		
+	0.5713	0.8409028		
+	0.5714	0.852104		
+	0.5715	0.845624		
+	0.5716	0.85648059		
+	0.5717	0.85347717		
+	0.5718	0.85028695		
+	0.5719	0.84745378		
+	0.572	0.86637144		
+	0.5721	0.85379985		
+	0.5722	0.86797191		
+	0.5723	0.87895375		
+	0.5724	0.87434247		
+	0.5725	0.87291644		
+	0.5726	0.88018685		
+	0.5727	0.88381779		
+	0.5728	0.89236302		
+	0.5729	0.88713007		
+	0.573	0.89244512		
+	0.5731	0.90960186		
+	0.5732	0.91872554		
+	0.5733	0.9221354		
+	0.5734	0.94084925		
+	0.5735	0.94188136		
+	0.5736	0.94674489		
+	0.5737	0.9433657		
+	0.5738	0.94490657		
+	0.5739	0.94555866		
+	0.574	0.94072211		
+	0.5741	0.92925042		
+	0.5742	0.93486296		
+	0.5743	0.93400332		
+	0.5744	0.91715145		
+	0.5745	0.91840333		
+	0.5746	0.91830568		
+	0.5747	0.91127331		
+	0.5748	0.91827283		
+	0.5749	0.90097093		
+	0.575	0.90625723		
+	0.5751	0.91045236		
+	0.5752	0.89673005		
+	0.5753	0.88952538		
+	0.5754	0.88704765		
+	0.5755	0.8957919		
+	0.5756	0.89190455		
+	0.5757	0.8886018		
+	0.5758	0.9017004		
+	0.5759	0.9060269		
+	0.576	0.91919961		
+	0.5761	0.91841865		
+	0.5762	0.94638422		
+	0.5763	0.94127501		
+	0.5764	0.93943249		
+	0.5765	0.95476783		
+	0.5766	0.94760784		
+	0.5767	0.94579092		
+	0.5768	0.94629795		
+	0.5769	0.93956304		
+	0.577	0.94127039		
+	0.5771	0.92555199		
+	0.5772	0.93047605		
+	0.5773	0.92921694		
+	0.5774	0.91883333		
+	0.5775	0.90833869		
+	0.5776	0.89853192		
+	0.5777	0.8968689		
+	0.5778	0.88240928		
+	0.5779	0.86866325		
+	0.578	0.8549186		
+	0.5781	0.84585623		
+	0.5782	0.84622973		
+	0.5783	0.84276873		
+	0.5784	0.82672369		
+	0.5785	0.81893007		
+	0.5786	0.82030453		
+	0.5787	0.81185015		
+	0.5788	0.81970823		
+	0.5789	0.82714561		
+	0.579	0.82731557		
+	0.5791	0.8373625		
+	0.5792	0.84104312		
+	0.5793	0.84113058		
+	0.5794	0.84402889		
+	0.5795	0.83994336		
+	0.5796	0.83881777		
+	0.5797	0.82590615		
+	0.5798	0.82253654		
+	0.5799	0.82075952		
+	0.58	0.83209364		
+	0.5801	0.81023765		
+	0.5802	0.80695081		
+	0.5803	0.81391806		
+	0.5804	0.81010026		
+	0.5805	0.79581576		
+	0.5806	0.80601462		
+	0.5807	0.78554708		
+	0.5808	0.79680624		
+	0.5809	0.7817549		
+	0.581	0.78603979		
+	0.5811	0.7911028		
+	0.5812	0.78925097		
+	0.5813	0.78671622		
+	0.5814	0.7789224		
+	0.5815	0.78289905		
+	0.5816	0.78219909		
+	0.5817	0.78401541		
+	0.5818	0.79996059		
+	0.5819	0.81784206		
+	0.582	0.82630709		
+	0.5821	0.81808997		
+	0.5822	0.83760935		
+	0.5823	0.8274617		
+	0.5824	0.82955265		
+	0.5825	0.82962558		
+	0.5826	0.83674092		
+	0.5827	0.82073131		
+	0.5828	0.81712759		
+	0.5829	0.81937771		
+	0.583	0.82776968		
+	0.5831	0.82385213		
+	0.5832	0.80778866		
+	0.5833	0.80543149		
+	0.5834	0.79882398		
+	0.5835	0.79870059		
+	0.5836	0.80272873		
+	0.5837	0.80147397		
+	0.5838	0.7977384		
+	0.5839	0.77952973		
+	0.584	0.78469019		
+	0.5841	0.78735191		
+	0.5842	0.77681149		
+	0.5843	0.77979794		
+	0.5844	0.78096568		
+	0.5845	0.78562497		
+	0.5846	0.7892996		
+	0.5847	0.80558161		
+	0.5848	0.80252658		
+	0.5849	0.82725194		
+	0.585	0.82967338		
+	0.5851	0.82786812		
+	0.5852	0.83737071		
+	0.5853	0.83269074		
+	0.5854	0.83931626		
+	0.5855	0.83522408		
+	0.5856	0.83586831		
+	0.5857	0.83395959		
+	0.5858	0.82479574		
+	0.5859	0.82672851		
+	0.586	0.81042542		
+	0.5861	0.82327202		
+	0.5862	0.81108076		
+	0.5863	0.79904662		
+	0.5864	0.80018144		
+	0.5865	0.80179806		
+	0.5866	0.78913938		
+	0.5867	0.79000253		
+	0.5868	0.80059693		
+	0.5869	0.78263702		
+	0.587	0.79040892		
+	0.5871	0.80154015		
+	0.5872	0.78936543		
+	0.5873	0.80306186		
+	0.5874	0.80827205		
+	0.5875	0.8075242		
+	0.5876	0.82618191		
+	0.5877	0.83323674		
+	0.5878	0.84441133		
+	0.5879	0.86073752		
+	0.588	0.87590277		
+	0.5881	0.88939112		
+	0.5882	0.90350079		
+	0.5883	0.89843039		
+	0.5884	0.90678796		
+	0.5885	0.91584844		
+	0.5886	0.9196198		
+	0.5887	0.91482868		
+	0.5888	0.91184233		
+	0.5889	0.922638		
+	0.589	0.90717362		
+	0.5891	0.91866208		
+	0.5892	0.91619572		
+	0.5893	0.89914818		
+	0.5894	0.89245143		
+	0.5895	0.8957388		
+	0.5896	0.89292838		
+	0.5897	0.9010228		
+	0.5898	0.88986018		
+	0.5899	0.89247504		
+	0.59	0.89625493		
+	0.5901	0.89093705		
+	0.5902	0.88518236		
+	0.5903	0.88560509		
+	0.5904	0.89751623		
+	0.5905	0.897039		
+	0.5906	0.91039289		
+	0.5907	0.91863718		
+	0.5908	0.9360235		
+	0.5909	0.94698163		
+	0.591	0.94957372		
+	0.5911	0.9519087		
+	0.5912	0.9434167		
+	0.5913	0.93993467		
+	0.5914	0.93182833		
+	0.5915	0.9499117		
+	0.5916	0.94112379		
+	0.5917	0.93047523		
+	0.5918	0.93575175		
+	0.5919	0.92701899		
+	0.592	0.91763091		
+	0.5921	0.92200601		
+	0.5922	0.9175218		
+	0.5923	0.91308918		
+	0.5924	0.90273254		
+	0.5925	0.9128235		
+	0.5926	0.90330115		
+	0.5927	0.90771241		
+	0.5928	0.89748319		
+	0.5929	0.90426727		
+	0.593	0.89477063		
+	0.5931	0.88547916		
+	0.5932	0.8955733		
+	0.5933	0.90107586		
+	0.5934	0.90187618		
+	0.5935	0.90944339		
+	0.5936	0.91992362		
+	0.5937	0.93663519		
+	0.5938	0.93434054		
+	0.5939	0.92946945		
+	0.594	0.93008119		
+	0.5941	0.90676443		
+	0.5942	0.90567615		
+	0.5943	0.89274094		
+	0.5944	0.89705634		
+	0.5945	0.89106266		
+	0.5946	0.86707543		
+	0.5947	0.86773201		
+	0.5948	0.85596792		
+	0.5949	0.84686575		
+	0.595	0.84444444		
+	0.5951	0.8273663		
+	0.5952	0.82146202		
+	0.5953	0.81571239		
+	0.5954	0.81767638		
+	0.5955	0.81210406		
+	0.5956	0.81093983		
+	0.5957	0.80182491		
+	0.5958	0.78819666		
+	0.5959	0.79941823		
+	0.596	0.78377518		
+	0.5961	0.77805756		
+	0.5962	0.78524726		
+	0.5963	0.78451955		
+	0.5964	0.79502202		
+	0.5965	0.80046588		
+	0.5966	0.82272855		
+	0.5967	0.81623155		
+	0.5968	0.83893742		
+	0.5969	0.82977267		
+	0.597	0.8299663		
+	0.5971	0.82103499		
+	0.5972	0.82683538		
+	0.5973	0.82941615		
+	0.5974	0.81792908		
+	0.5975	0.82447905		
+	0.5976	0.82417979		
+	0.5977	0.80696706		
+	0.5978	0.81664843		
+	0.5979	0.81447052		
+	0.598	0.80789273		
+	0.5981	0.81074836		
+	0.5982	0.80599141		
+	0.5983	0.80208847		
+	0.5984	0.79835902		
+	0.5985	0.78640155		
+	0.5986	0.79531024		
+	0.5987	0.79008969		
+	0.5988	0.78975914		
+	0.5989	0.78987768		
+	0.599	0.78935276		
+	0.5991	0.77499228		
+	0.5992	0.79087191		
+	0.5993	0.79552231		
+	0.5994	0.80492092		
+	0.5995	0.81013644		
+	0.5996	0.81831584		
+	0.5997	0.82660142		
+	0.5998	0.83711736		
+	0.5999	0.84195454		
+	0.6	0.84129557		
+	0.6001	0.82773139		
+	0.6002	0.83086553		
+	0.6003	0.83027381		
+	0.6004	0.81599701		
+	0.6005	0.83057624		
+	0.6006	0.82039018		
+	0.6007	0.80708343		
+	0.6008	0.80750091		
+	0.6009	0.81263984		
+	0.601	0.79700408		
+	0.6011	0.79232307		
+	0.6012	0.79528282		
+	0.6013	0.80338789		
+	0.6014	0.80024613		
+	0.6015	0.78722487		
+	0.6016	0.78309662		
+	0.6017	0.78164248		
+	0.6018	0.79380176		
+	0.6019	0.7777953		
+	0.602	0.77699689		
+	0.6021	0.78567614		
+	0.6022	0.79212348		
+	0.6023	0.80954493		
+	0.6024	0.82120239		
+	0.6025	0.81723548		
+	0.6026	0.84112549		
+	0.6027	0.84317889		
+	0.6028	0.83099505		
+	0.6029	0.82744299		
+	0.603	0.84435063		
+	0.6031	0.8241198		
+	0.6032	0.8378344		
+	0.6033	0.83594128		
+	0.6034	0.83971075		
+	0.6035	0.83509409		
+	0.6036	0.83429102		
+	0.6037	0.8307441		
+	0.6038	0.84092299		
+	0.6039	0.82672256		
+	0.604	0.84267506		
+	0.6041	0.84572613		
+	0.6042	0.84211896		
+	0.6043	0.84799195		
+	0.6044	0.84713283		
+	0.6045	0.8465939		
+	0.6046	0.85953612		
+	0.6047	0.8566473		
+	0.6048	0.85635837		
+	0.6049	0.86831336		
+	0.605	0.87131034		
+	0.6051	0.89195861		
+	0.6052	0.91118375		
+	0.6053	0.91861501		
+	0.6054	0.92496087		
+	0.6055	0.94349549		
+	0.6056	0.94448346		
+	0.6057	0.933382		
+	0.6058	0.94160876		
+	0.6059	0.94148744		
+	0.606	0.93407094		
+	0.6061	0.94323384		
+	0.6062	0.93809135		
+	0.6063	0.93733881		
+	0.6064	0.93064423		
+	0.6065	0.93702734		
+	0.6066	0.92021802		
+	0.6067	0.93161043		
+	0.6068	0.91885385		
+	0.6069	0.91018068		
+	0.607	0.91449286		
+	0.6071	0.91482123		
+	0.6072	0.90649574		
+	0.6073	0.89899014		
+	0.6074	0.90777905		
+	0.6075	0.90493432		
+	0.6076	0.90512127		
+	0.6077	0.89203493		
+	0.6078	0.89223723		
+	0.6079	0.90228454		
+	0.608	0.90613608		
+	0.6081	0.91305106		
+	0.6082	0.92945492		
+	0.6083	0.94069958		
+	0.6084	0.94341866		
+	0.6085	0.94535092		
+	0.6086	0.95370934		
+	0.6087	0.94554464		
+	0.6088	0.94791767		
+	0.6089	0.95290051		
+	0.609	0.94254185		
+	0.6091	0.95227223		
+	0.6092	0.93944724		
+	0.6093	0.94303082		
+	0.6094	0.93783338		
+	0.6095	0.93358026		
+	0.6096	0.91890142		
+	0.6097	0.92762197		
+	0.6098	0.92062319		
+	0.6099	0.91967161		
+	0.61	0.91190226		
+	0.6101	0.89880123		
+	0.6102	0.89566245		
+	0.6103	0.87621791		
+	0.6104	0.86876522		
+	0.6105	0.85648295		
+	0.6106	0.8636001		
+	0.6107	0.85358745		
+	0.6108	0.85153572		
+	0.6109	0.83532873		
+	0.611	0.8503959		
+	0.6111	0.85943917		
+	0.6112	0.85986303		
+	0.6113	0.85780497		
+	0.6114	0.86503571		
+	0.6115	0.8546113		
+	0.6116	0.85074613		
+	0.6117	0.86082668		
+	0.6118	0.85859672		
+	0.6119	0.85108928		
+	0.612	0.83706185		
+	0.6121	0.84430256		
+	0.6122	0.83998275		
+	0.6123	0.81957618		
+	0.6124	0.81274101		
+	0.6125	0.82100726		
+	0.6126	0.81583526		
+	0.6127	0.8001195		
+	0.6128	0.79877598		
+	0.6129	0.79586605		
+	0.613	0.79324677		
+	0.6131	0.79803589		
+	0.6132	0.7834458		
+	0.6133	0.79455819		
+	0.6134	0.79400059		
+	0.6135	0.78533231		
+	0.6136	0.79446168		
+	0.6137	0.78150755		
+	0.6138	0.79819021		
+	0.6139	0.79516449		
+	0.614	0.80761066		
+	0.6141	0.82414324		
+	0.6142	0.82313636		
+	0.6143	0.82813183		
+	0.6144	0.84267066		
+	0.6145	0.82887653		
+	0.6146	0.83524508		
+	0.6147	0.84370264		
+	0.6148	0.83726332		
+	0.6149	0.83359961		
+	0.615	0.83181186		
+	0.6151	0.82238594		
+	0.6152	0.81591592		
+	0.6153	0.82748867		
+	0.6154	0.81119041		
+	0.6155	0.81219668		
+	0.6156	0.80572949		
+	0.6157	0.81232156		
+	0.6158	0.79627592		
+	0.6159	0.79208019		
+	0.616	0.78601357		
+	0.6161	0.79475875		
+	0.6162	0.79966245		
+	0.6163	0.79310699		
+	0.6164	0.78457592		
+	0.6165	0.78871325		
+	0.6166	0.78148875		
+	0.6167	0.7855076		
+	0.6168	0.79789597		
+	0.6169	0.79850877		
+	0.617	0.81903007		
+	0.6171	0.82784838		
+	0.6172	0.8384479		
+	0.6173	0.84417324		
+	0.6174	0.84906899		
+	0.6175	0.84805206		
+	0.6176	0.82901264		
+	0.6177	0.83869007		
+	0.6178	0.83309731		
+	0.6179	0.84265214		
+	0.618	0.83748584		
+	0.6181	0.82835477		
+	0.6182	0.83216018		
+	0.6183	0.81241781		
+	0.6184	0.82195349		
+	0.6185	0.81350568		
+	0.6186	0.80979676		
+	0.6187	0.79889737		
+	0.6188	0.79589717		
+	0.6189	0.80364759		
+	0.619	0.79477094		
+	0.6191	0.78529662		
+	0.6192	0.79149738		
+	0.6193	0.80145946		
+	0.6194	0.78537716		
+	0.6195	0.79046433		
+	0.6196	0.80071426		
+	0.6197	0.81624161		
+	0.6198	0.81402		
+	0.6199	0.82667185		
+	0.62	0.85558448		
+	0.6201	0.86548138		
+	0.6202	0.86560622		
+	0.6203	0.87802826		
+	0.6204	0.89145709		
+	0.6205	0.891366		
+	0.6206	0.88288217		
+	0.6207	0.9020952		
+	0.6208	0.89951051		
+	0.6209	0.90882624		
+	0.621	0.91559298		
+	0.6211	0.91752699		
+	0.6212	0.90418605		
+	0.6213	0.91111004		
+	0.6214	0.9133172		
+	0.6215	0.90749616		
+	0.6216	0.90106808		
+	0.6217	0.90843744		
+	0.6218	0.90457842		
+	0.6219	0.90413754		
+	0.622	0.8925593		
+	0.6221	0.89520479		
+	0.6222	0.88895577		
+	0.6223	0.90493299		
+	0.6224	0.89484859		
+	0.6225	0.90553761		
+	0.6226	0.90677041		
+	0.6227	0.91689765		
+	0.6228	0.92081362		
+	0.6229	0.92954043		
+	0.623	0.95184175		
+	0.6231	0.95227564		
+	0.6232	0.95176299		
+	0.6233	0.95887129		
+	0.6234	0.95899416		
+	0.6235	0.94608672		
+	0.6236	0.95434931		
+	0.6237	0.95133819		
+	0.6238	0.94018998		
+	0.6239	0.95063694		
+	0.624	0.93426506		
+	0.6241	0.94622637		
+	0.6242	0.93589634		
+	0.6243	0.92010295		
+	0.6244	0.92256611		
+	0.6245	0.91688965		
+	0.6246	0.91046114		
+	0.6247	0.91061022		
+	0.6248	0.92114658		
+	0.6249	0.9060722		
+	0.625	0.90592853		
+	0.6251	0.9049429		
+	0.6252	0.91284244		
+	0.6253	0.9001406		
+	0.6254	0.89801083		
+	0.6255	0.91445753		
+	0.6256	0.91338351		
+	0.6257	0.93281809		
+	0.6258	0.93320569		
+	0.6259	0.95606865		
+	0.626	0.94551637		
+	0.6261	0.95503804		
+	0.6262	0.96426419		
+	0.6263	0.95792169		
+	0.6264	0.9409664		
+	0.6265	0.93291867		
+	0.6266	0.93243406		
+	0.6267	0.91944867		
+	0.6268	0.90009525		
+	0.6269	0.90102278		
+	0.627	0.89724889		
+	0.6271	0.87392323		
+	0.6272	0.87612148		
+	0.6273	0.86032245		
+	0.6274	0.85359568		
+	0.6275	0.84058139		
+	0.6276	0.83905172		
+	0.6277	0.82282239		
+	0.6278	0.82806154		
+	0.6279	0.82578897		
+	0.628	0.81349487		
+	0.6281	0.81478567		
+	0.6282	0.80476666		
+	0.6283	0.80155819		
+	0.6284	0.80574553		
+	0.6285	0.80605541		
+	0.6286	0.8146852		
+	0.6287	0.82231186		
+	0.6288	0.83900007		
+	0.6289	0.83312395		
+	0.629	0.8365502		
+	0.6291	0.83562337		
+	0.6292	0.84764161		
+	0.6293	0.84412489		
+	0.6294	0.84573181		
+	0.6295	0.83149066		
+	0.6296	0.83356381		
+	0.6297	0.82684289		
+	0.6298	0.82423956		
+	0.6299	0.82838677		
+	0.63	0.82148192		
+	0.6301	0.82868882		
+	0.6302	0.8085623		
+	0.6303	0.80952001		
+	0.6304	0.80106067		
+	0.6305	0.80960911		
+	0.6306	0.80419174		
+	0.6307	0.79925191		
+	0.6308	0.79363292		
+	0.6309	0.80507865		
+	0.631	0.80275634		
+	0.6311	0.78738876		
+	0.6312	0.78464954		
+	0.6313	0.79409105		
+	0.6314	0.80162228		
+	0.6315	0.81259424		
+	0.6316	0.8286079		
+	0.6317	0.83695725		
+	0.6318	0.83358353		
+	0.6319	0.84593165		
+	0.632	0.843972		
+	0.6321	0.85112908		
+	0.6322	0.84842026		
+	0.6323	0.84369934		
+	0.6324	0.84041935		
+	0.6325	0.84509795		
+	0.6326	0.83348837		
+	0.6327	0.84113492		
+	0.6328	0.83125105		
+	0.6329	0.81972644		
+	0.633	0.81870583		
+	0.6331	0.81112569		
+	0.6332	0.82316097		
+	0.6333	0.80582078		
+	0.6334	0.8114868		
+	0.6335	0.80269081		
+	0.6336	0.81227028		
+	0.6337	0.79973702		
+	0.6338	0.79207361		
+	0.6339	0.78884229		
+	0.634	0.80076796		
+	0.6341	0.79344685		
+	0.6342	0.79064491		
+	0.6343	0.79588301		
+	0.6344	0.82191982		
+	0.6345	0.82521188		
+	0.6346	0.83052539		
+	0.6347	0.8370614		
+	0.6348	0.83823964		
+	0.6349	0.84116221		
+	0.635	0.84348843		
+	0.6351	0.85577986		
+	0.6352	0.85221377		
+	0.6353	0.85145685		
+	0.6354	0.83557899		
+	0.6355	0.84344894		
+	0.6356	0.8370788		
+	0.6357	0.84121616		
+	0.6358	0.84587045		
+	0.6359	0.83575635		
+	0.636	0.82798927		
+	0.6361	0.84348298		
+	0.6362	0.84351933		
+	0.6363	0.82910071		
+	0.6364	0.83908132		
+	0.6365	0.82931913		
+	0.6366	0.83535199		
+	0.6367	0.84345636		
+	0.6368	0.84390175		
+	0.6369	0.8479152		
+	0.637	0.86015038		
+	0.6371	0.87285491		
+	0.6372	0.87584316		
+	0.6373	0.89494832		
+	0.6374	0.91174045		
+	0.6375	0.92111923		
+	0.6376	0.93258103		
+	0.6377	0.95464985		
+	0.6378	0.95141881		
+	0.6379	0.94645566		
+	0.638	0.94722444		
+	0.6381	0.95212567		
+	0.6382	0.94835673		
+	0.6383	0.95566299		
+	0.6384	0.94648232		
+	0.6385	0.94536487		
+	0.6386	0.9463043		
+	0.6387	0.94674382		
+	0.6388	0.93242381		
+	0.6389	0.92516214		
+	0.639	0.93544552		
+	0.6391	0.936855		
+	0.6392	0.9263223		
+	0.6393	0.92732294		
+	0.6394	0.92657473		
+	0.6395	0.91179009		
+	0.6396	0.91357122		
+	0.6397	0.91310783		
+	0.6398	0.90421218		
+	0.6399	0.91871328		
+	0.64	0.9142994		
+	0.6401	0.91675514		
+	0.6402	0.92913072		
+	0.6403	0.93079356		
+	0.6404	0.94083384		
+	0.6405	0.96423781		
+	0.6406	0.95410125		
+	0.6407	0.95986992		
+	0.6408	0.96689566		
+	0.6409	0.96165809		
+	0.641	0.95915459		
+	0.6411	0.96203497		
+	0.6412	0.95694341		
+	0.6413	0.96019515		
+	0.6414	0.95402425		
+	0.6415	0.95218962		
+	0.6416	0.94971403		
+	0.6417	0.94931154		
+	0.6418	0.94198741		
+	0.6419	0.93055009		
+	0.642	0.92518823		
+	0.6421	0.9363201		
+	0.6422	0.91832876		
+	0.6423	0.92834491		
+	0.6424	0.91416792		
+	0.6425	0.9239145		
+	0.6426	0.90722637		
+	0.6427	0.90120351		
+	0.6428	0.89726375		
+	0.6429	0.89815878		
+	0.643	0.88578232		
+	0.6431	0.89201936		
+	0.6432	0.89532553		
+	0.6433	0.88376953		
+	0.6434	0.90507745		
+	0.6435	0.90646942		
+	0.6436	0.89292499		
+	0.6437	0.89501031		
+	0.6438	0.8848365		
+	0.6439	0.87454936		
+	0.644	0.86995193		
+	0.6441	0.86786617		
+	0.6442	0.86200075		
+	0.6443	0.86711506		
+	0.6444	0.86268248		
+	0.6445	0.84967687		
+	0.6446	0.85126996		
+	0.6447	0.82975988		
+	0.6448	0.82447105		
+	0.6449	0.83455011		
+	0.645	0.82944665		
+	0.6451	0.81718067		
+	0.6452	0.81291801		
+	0.6453	0.80480721		
+	0.6454	0.81756126		
+	0.6455	0.8066901		
+	0.6456	0.80490664		
+	0.6457	0.80562071		
+	0.6458	0.80505194		
+	0.6459	0.79518855		
+	0.646	0.81643221		
+	0.6461	0.81028701		
+	0.6462	0.82246194		
+	0.6463	0.83389542		
+	0.6464	0.83818054		
+	0.6465	0.84629713		
+	0.6466	0.84623385		
+	0.6467	0.85217769		
+	0.6468	0.85708201		
+	0.6469	0.8567446		
+	0.647	0.84397		
+	0.6471	0.8411962		
+	0.6472	0.84360427		
+	0.6473	0.85164803		
+	0.6474	0.83758627		
+	0.6475	0.83889725		
+	0.6476	0.83908113		
+	0.6477	0.82115717		
+	0.6478	0.83319016		
+	0.6479	0.81550897		
+	0.648	0.81442246		
+	0.6481	0.8239775		
+	0.6482	0.8133857		
+	0.6483	0.81338665		
+	0.6484	0.81440198		
+	0.6485	0.8047117		
+	0.6486	0.79734789		
+	0.6487	0.80509079		
+	0.6488	0.80299029		
+	0.6489	0.80896904		
+	0.649	0.82178852		
+	0.6491	0.82720408		
+	0.6492	0.84974371		
+	0.6493	0.85439179		
+	0.6494	0.85985144		
+	0.6495	0.8588883		
+	0.6496	0.85178063		
+	0.6497	0.86209488		
+	0.6498	0.8608868		
+	0.6499	0.8517422		
+	0.65	0.85779735		
+	0.6501	0.85031934		
+	0.6502	0.85617243		
+	0.6503	0.85073044		
+	0.6504	0.83217489		
+	0.6505	0.82843373		
+	0.6506	0.8378772		
+	0.6507	0.83464655		
+	0.6508	0.83426104		
+	0.6509	0.81902767		
+	0.651	0.81062353		
+	0.6511	0.8159021		
+	0.6512	0.81739442		
+	0.6513	0.80440405		
+	0.6514	0.80880588		
+	0.6515	0.81242047		
+	0.6516	0.80987871		
+	0.6517	0.8113753		
+	0.6518	0.81648442		
+	0.6519	0.81333971		
+	0.652	0.83829638		
+	0.6521	0.84483674		
+	0.6522	0.85255437		
+	0.6523	0.87729349		
+	0.6524	0.8817591		
+	0.6525	0.87840356		
+	0.6526	0.88351175		
+	0.6527	0.8903801		
+	0.6528	0.88253059		
+	0.6529	0.88463214		
+	0.653	0.88774994		
+	0.6531	0.90103387		
+	0.6532	0.90835913		
+	0.6533	0.90007209		
+	0.6534	0.90472641		
+	0.6535	0.90673724		
+	0.6536	0.9096422		
+	0.6537	0.90912505		
+	0.6538	0.9091828		
+	0.6539	0.91051629		
+	0.654	0.90632986		
+	0.6541	0.91126102		
+	0.6542	0.91306587		
+	0.6543	0.91228009		
+	0.6544	0.9064441		
+	0.6545	0.91739161		
+	0.6546	0.90852652		
+	0.6547	0.91344889		
+	0.6548	0.92868212		
+	0.6549	0.9440238		
+	0.655	0.9517207		
+	0.6551	0.96116394		
+	0.6552	0.97383641		
+	0.6553	0.97129412		
+	0.6554	0.97513716		
+	0.6555	0.96234418		
+	0.6556	0.97091392		
+	0.6557	0.97629268		
+	0.6558	0.97334016		
+	0.6559	0.97372312		
+	0.656	0.96153473		
+	0.6561	0.96594671		
+	0.6562	0.95737428		
+	0.6563	0.9520895		
+	0.6564	0.95000823		
+	0.6565	0.9434413		
+	0.6566	0.94297824		
+	0.6567	0.93734405		
+	0.6568	0.93753783		
+	0.6569	0.94366727		
+	0.657	0.93132954		
+	0.6571	0.92386913		
+	0.6572	0.93596236		
+	0.6573	0.93003017		
+	0.6574	0.92627937		
+	0.6575	0.93370745		
+	0.6576	0.92046504		
+	0.6577	0.92856145		
+	0.6578	0.94705751		
+	0.6579	0.9589636		
+	0.658	0.95634429		
+	0.6581	0.97937164		
+	0.6582	0.97426525		
+	0.6583	0.98534503		
+	0.6584	0.98293048		
+	0.6585	0.98271701		
+	0.6586	0.97783229		
+	0.6587	0.9672525		
+	0.6588	0.96268349		
+	0.6589	0.96340585		
+	0.659	0.95222344		
+	0.6591	0.94115707		
+	0.6592	0.9415522		
+	0.6593	0.91604185		
+	0.6594	0.91198344		
+	0.6595	0.90721602		
+	0.6596	0.88606696		
+	0.6597	0.88428203		
+	0.6598	0.88320705		
+	0.6599	0.85750943		
+	0.66	0.85824987		
+	0.6601	0.84881439		
+	0.6602	0.84584002		
+	0.6603	0.83812015		
+	0.6604	0.83481894		
+	0.6605	0.83332751		
+	0.6606	0.84601851		
+	0.6607	0.83434165		
+	0.6608	0.84161762		
+	0.6609	0.85594326		
+	0.661	0.86909392		
+	0.6611	0.86657289		
+	0.6612	0.86468439		
+	0.6613	0.86276322		
+	0.6614	0.86111213		
+	0.6615	0.86919363		
+	0.6616	0.86244006		
+	0.6617	0.85363047		
+	0.6618	0.84692666		
+	0.6619	0.84796738		
+	0.662	0.84497345		
+	0.6621	0.84588128		
+	0.6622	0.84448223		
+	0.6623	0.83814255		
+	0.6624	0.82685237		
+	0.6625	0.83169568		
+	0.6626	0.82258528		
+	0.6627	0.82380052		
+	0.6628	0.81878964		
+	0.6629	0.80995608		
+	0.663	0.80846167		
+	0.6631	0.82301801		
+	0.6632	0.82003136		
+	0.6633	0.81738909		
+	0.6634	0.82045669		
+	0.6635	0.81683272		
+	0.6636	0.82772046		
+	0.6637	0.83783069		
+	0.6638	0.84689569		
+	0.6639	0.8624409		
+	0.664	0.85821555		
+	0.6641	0.86282865		
+	0.6642	0.87130296		
+	0.6643	0.86381138		
+	0.6644	0.87205118		
+	0.6645	0.86592952		
+	0.6646	0.85319039		
+	0.6647	0.85127367		
+	0.6648	0.85841659		
+	0.6649	0.86213617		
+	0.665	0.85944882		
+	0.6651	0.84228233		
+	0.6652	0.84299072		
+	0.6653	0.83536785		
+	0.6654	0.83292506		
+	0.6655	0.82375832		
+	0.6656	0.82821455		
+	0.6657	0.82798941		
+	0.6658	0.82842607		
+	0.6659	0.81685342		
+	0.666	0.8109982		
+	0.6661	0.82650172		
+	0.6662	0.81361377		
+	0.6663	0.82396956		
+	0.6664	0.82564871		
+	0.6665	0.8248307		
+	0.6666	0.83513943		
+	0.6667	0.8479554		
+	0.6668	0.85112986		
+	0.6669	0.8606517		
+	0.667	0.8732075		
+	0.6671	0.86350276		
+	0.6672	0.86621244		
+	0.6673	0.86626314		
+	0.6674	0.85759965		
+	0.6675	0.87417953		
+	0.6676	0.85467684		
+	0.6677	0.85481755		
+	0.6678	0.85759459		
+	0.6679	0.84909836		
+	0.668	0.84195231		
+	0.6681	0.85549067		
+	0.6682	0.84521891		
+	0.6683	0.84120734		
+	0.6684	0.83724665		
+	0.6685	0.83600006		
+	0.6686	0.8317584		
+	0.6687	0.83799307		
+	0.6688	0.84188848		
+	0.6689	0.84146913		
+	0.669	0.85751094		
+	0.6691	0.84554964		
+	0.6692	0.8669228		
+	0.6693	0.86026351		
+	0.6694	0.87091042		
+	0.6695	0.88525715		
+	0.6696	0.90704341		
+	0.6697	0.91777736		
+	0.6698	0.9344277		
+	0.6699	0.94812572		
+	0.67	0.95089748		
+	0.6701	0.95629639		
+	0.6702	0.96715376		
+	0.6703	0.97680603		
+	0.6704	0.97415091		
+	0.6705	0.97044932		
+	0.6706	0.96413144		
+	0.6707	0.96670468		
+	0.6708	0.966404		
+	0.6709	0.95404491		
+	0.671	0.960568		
+	0.6711	0.94479902		
+	0.6712	0.94583779		
+	0.6713	0.95177333		
+	0.6714	0.94599141		
+	0.6715	0.94906037		
+	0.6716	0.94716822		
+	0.6717	0.92710164		
+	0.6718	0.93708167		
+	0.6719	0.94127704		
+	0.672	0.93993158		
+	0.6721	0.94237416		
+	0.6722	0.9312371		
+	0.6723	0.95033363		
+	0.6724	0.93903518		
+	0.6725	0.95950207		
+	0.6726	0.9673598		
+	0.6727	0.98849624		
+	0.6728	0.98354942		
+	0.6729	0.99227054		
+	0.673	0.9818896		
+	0.6731	0.99510329		
+	0.6732	0.98652402		
+	0.6733	0.99141497		
+	0.6734	0.97496705		
+	0.6735	0.97139521		
+	0.6736	0.98346422		
+	0.6737	0.97753398		
+	0.6738	0.97611032		
+	0.6739	0.97512483		
+	0.674	0.9687931		
+	0.6741	0.95904037		
+	0.6742	0.94941395		
+	0.6743	0.94728795		
+	0.6744	0.94726044		
+	0.6745	0.94681876		
+	0.6746	0.94176077		
+	0.6747	0.94358447		
+	0.6748	0.9392864		
+	0.6749	0.93875699		
+	0.675	0.94030267		
+	0.6751	0.93366757		
+	0.6752	0.94432608		
+	0.6753	0.93186649		
+	0.6754	0.9523246		
+	0.6755	0.9524082		
+	0.6756	0.95017353		
+	0.6757	0.94800327		
+	0.6758	0.93830907		
+	0.6759	0.93527406		
+	0.676	0.92141617		
+	0.6761	0.92737382		
+	0.6762	0.91777813		
+	0.6763	0.90124667		
+	0.6764	0.90326482		
+	0.6765	0.9069978		
+	0.6766	0.89364524		
+	0.6767	0.87625222		
+	0.6768	0.87655775		
+	0.6769	0.86179779		
+	0.677	0.85412045		
+	0.6771	0.85601809		
+	0.6772	0.85458608		
+	0.6773	0.83922378		
+	0.6774	0.84932031		
+	0.6775	0.84589982		
+	0.6776	0.82679014		
+	0.6777	0.82148249		
+	0.6778	0.81857201		
+	0.6779	0.82048686		
+	0.678	0.8173201		
+	0.6781	0.82429042		
+	0.6782	0.83009448		
+	0.6783	0.83586015		
+	0.6784	0.85939949		
+	0.6785	0.86280416		
+	0.6786	0.87152836		
+	0.6787	0.87801744		
+	0.6788	0.87002669		
+	0.6789	0.8711758		
+	0.679	0.87670364		
+	0.6791	0.87999567		
+	0.6792	0.86299583		
+	0.6793	0.87779556		
+	0.6794	0.87404834		
+	0.6795	0.86858823		
+	0.6796	0.860897		
+	0.6797	0.8526647		
+	0.6798	0.84364839		
+	0.6799	0.8391047		
+	0.68	0.84074975		
+	0.6801	0.83894592		
+	0.6802	0.84430268		
+	0.6803	0.83196036		
+	0.6804	0.83307717		
+	0.6805	0.82197821		
+	0.6806	0.83151256		
+	0.6807	0.82678286		
+	0.6808	0.82212658		
+	0.6809	0.8175062		
+	0.681	0.83566819		
+	0.6811	0.83779832		
+	0.6812	0.85188568		
+	0.6813	0.85676847		
+	0.6814	0.87378037		
+	0.6815	0.87519859		
+	0.6816	0.88265901		
+	0.6817	0.8861409		
+	0.6818	0.88171274		
+	0.6819	0.8824877		
+	0.682	0.86817212		
+	0.6821	0.88487065		
+	0.6822	0.8675825		
+	0.6823	0.86235579		
+	0.6824	0.86446047		
+	0.6825	0.85949191		
+	0.6826	0.85157256		
+	0.6827	0.85962103		
+	0.6828	0.84924438		
+	0.6829	0.85412792		
+	0.683	0.85148936		
+	0.6831	0.84825694		
+	0.6832	0.84139964		
+	0.6833	0.82984258		
+	0.6834	0.83123219		
+	0.6835	0.83215049		
+	0.6836	0.83906411		
+	0.6837	0.8354707		
+	0.6838	0.83750054		
+	0.6839	0.83928019		
+	0.684	0.83027434		
+	0.6841	0.85384657		
+	0.6842	0.8474574		
+	0.6843	0.86793967		
+	0.6844	0.87753898		
+	0.6845	0.88622658		
+	0.6846	0.88560355		
+	0.6847	0.88538654		
+	0.6848	0.89044106		
+	0.6849	0.89557426		
+	0.685	0.90128155		
+	0.6851	0.89024438		
+	0.6852	0.89846486		
+	0.6853	0.90410127		
+	0.6854	0.90601104		
+	0.6855	0.89742134		
+	0.6856	0.89541081		
+	0.6857	0.90508056		
+	0.6858	0.90274594		
+	0.6859	0.91334256		
+	0.686	0.90989616		
+	0.6861	0.92380152		
+	0.6862	0.92066871		
+	0.6863	0.93255065		
+	0.6864	0.91943353		
+	0.6865	0.92809039		
+	0.6866	0.93438373		
+	0.6867	0.92600986		
+	0.6868	0.92974548		
+	0.6869	0.94424664		
+	0.687	0.94405579		
+	0.6871	0.96188842		
+	0.6872	0.96226748		
+	0.6873	0.97806315		
+	0.6874	0.98384589		
+	0.6875	0.99203135		
+	0.6876	0.99512737		
+	0.6877	0.98433298		
+	0.6878	0.99089068		
+	0.6879	0.99486297		
+	0.688	0.99206968		
+	0.6881	0.99094527		
+	0.6882	0.98393808		
+	0.6883	0.97923633		
+	0.6884	0.97888026		
+	0.6885	0.9710276		
+	0.6886	0.97051924		
+	0.6887	0.96367091		
+	0.6888	0.96023395		
+	0.6889	0.96203265		
+	0.689	0.96061749		
+	0.6891	0.94991193		
+	0.6892	0.95806211		
+	0.6893	0.94953506		
+	0.6894	0.94207256		
+	0.6895	0.93981677		
+	0.6896	0.95314651		
+	0.6897	0.9482944		
+	0.6898	0.94563741		
+	0.6899	0.94787349		
+	0.69	0.96942101		
+	0.6901	0.97012193		
+	0.6902	0.97870378		
+	0.6903	0.99889016		
+	0.6904	1.0017916		
+	0.6905	1.003478		
+	0.6906	1.0063236		
+	0.6907	1.0010132		
+	0.6908	0.99972777		
+	0.6909	0.98608093		
+	0.691	0.99173465		
+	0.6911	0.9886147		
+	0.6912	0.99060651		
+	0.6913	0.98411783		
+	0.6914	0.96832459		
+	0.6915	0.9777239		
+	0.6916	0.96329205		
+	0.6917	0.95466983		
+	0.6918	0.9378912		
+	0.6919	0.93810214		
+	0.692	0.9162636		
+	0.6921	0.91086204		
+	0.6922	0.907037		
+	0.6923	0.89183522		
+	0.6924	0.88649622		
+	0.6925	0.88346055		
+	0.6926	0.87512403		
+	0.6927	0.86780788		
+	0.6928	0.8787568		
+	0.6929	0.88848577		
+	0.693	0.89320936		
+	0.6931	0.89788123		
+	0.6932	0.90227047		
+	0.6933	0.89983295		
+	0.6934	0.89907809		
+	0.6935	0.88889972		
+	0.6936	0.89183189		
+	0.6937	0.89531476		
+	0.6938	0.89128206		
+	0.6939	0.87930609		
+	0.694	0.8844303		
+	0.6941	0.87360307		
+	0.6942	0.86515164		
+	0.6943	0.85841551		
+	0.6944	0.85633087		
+	0.6945	0.85296134		
+	0.6946	0.85568228		
+	0.6947	0.85960731		
+	0.6948	0.85227609		
+	0.6949	0.84898182		
+	0.695	0.84421872		
+	0.6951	0.84066911		
+	0.6952	0.82871426		
+	0.6953	0.83883531		
+	0.6954	0.83871365		
+	0.6955	0.84216008		
+	0.6956	0.83498259		
+	0.6957	0.85210624		
+	0.6958	0.84528653		
+	0.6959	0.86721043		
+	0.696	0.86650997		
+	0.6961	0.88635607		
+	0.6962	0.8830679		
+	0.6963	0.89518737		
+	0.6964	0.88527913		
+	0.6965	0.88683378		
+	0.6966	0.87771952		
+	0.6967	0.88265588		
+	0.6968	0.89013255		
+	0.6969	0.88888052		
+	0.697	0.8721328		
+	0.6971	0.8656887		
+	0.6972	0.87474777		
+	0.6973	0.85697947		
+	0.6974	0.87114525		
+	0.6975	0.86297574		
+	0.6976	0.84840939		
+	0.6977	0.85639484		
+	0.6978	0.84375932		
+	0.6979	0.84408953		
+	0.698	0.83548758		
+	0.6981	0.8473207		
+	0.6982	0.83789468		
+	0.6983	0.8318948		
+	0.6984	0.83505724		
+	0.6985	0.83367617		
+	0.6986	0.85334188		
+	0.6987	0.84349658		
+	0.6988	0.8680884		
+	0.6989	0.88178853		
+	0.699	0.8812047		
+	0.6991	0.8832383		
+	0.6992	0.89217947		
+	0.6993	0.89243823		
+	0.6994	0.89461867		
+	0.6995	0.89359511		
+	0.6996	0.88043103		
+	0.6997	0.88690688		
+	0.6998	0.89324892		
+	0.6999	0.89085897		
+	0.7	0.87865077		
+	0.7001	0.86482958		
+	0.7002	0.86272835		
+	0.7003	0.86678586		
+	0.7004	0.8581388		
+	0.7005	0.86580462		
+	0.7006	0.84947506		
+	0.7007	0.85762858		
+	0.7008	0.84757149		
+	0.7009	0.85674202		
+	0.701	0.84463318		
+	0.7011	0.84272628		
+	0.7012	0.85905234		
+	0.7013	0.85506904		
+	0.7014	0.85240329		
+	0.7015	0.86934619		
+	0.7016	0.88959318		
+	0.7017	0.89299048		
+	0.7018	0.90831196		
+	0.7019	0.92024734		
+	0.702	0.93305953		
+	0.7021	0.94087089		
+	0.7022	0.95016955		
+	0.7023	0.96926794		
+	0.7024	0.95576993		
+	0.7025	0.97083296		
+	0.7026	0.98253707		
+	0.7027	0.97799992		
+	0.7028	0.97248622		
+	0.7029	0.98134357		
+	0.703	0.98282062		
+	0.7031	0.96376802		
+	0.7032	0.97097568		
+	0.7033	0.95859887		
+	0.7034	0.95558751		
+	0.7035	0.96547576		
+	0.7036	0.95927728		
+	0.7037	0.94852512		
+	0.7038	0.95007643		
+	0.7039	0.9533694		
+	0.704	0.95928036		
+	0.7041	0.95417842		
+	0.7042	0.95018082		
+	0.7043	0.95781829		
+	0.7044	0.95037012		
+	0.7045	0.95809145		
+	0.7046	0.97200107		
+	0.7047	0.98371747		
+	0.7048	0.99131735		
+	0.7049	0.99599272		
+	0.705	1.0147073		
+	0.7051	1.01097		
+	0.7052	0.9978337		
+	0.7053	1.0084851		
+	0.7054	1.0002697		
+	0.7055	1.007258		
+	0.7056	1.0090583		
+	0.7057	0.993749		
+	0.7058	0.98747468		
+	0.7059	0.98540507		
+	0.706	0.97917858		
+	0.7061	0.9903156		
+	0.7062	0.97376959		
+	0.7063	0.96714866		
+	0.7064	0.98031179		
+	0.7065	0.963221		
+	0.7066	0.97486074		
+	0.7067	0.96563999		
+	0.7068	0.95805313		
+	0.7069	0.96882806		
+	0.707	0.95929916		
+	0.7071	0.96434781		
+	0.7072	0.96273904		
+	0.7073	0.96258265		
+	0.7074	0.95623399		
+	0.7075	0.96949076		
+	0.7076	0.97135427		
+	0.7077	0.99318898		
+	0.7078	0.98853381		
+	0.7079	0.99754092		
+	0.708	1.0017098		
+	0.7081	0.9930251		
+	0.7082	0.97110318		
+	0.7083	0.97593331		
+	0.7084	0.95958207		
+	0.7085	0.95197125		
+	0.7086	0.93758122		
+	0.7087	0.92920673		
+	0.7088	0.9215455		
+	0.7089	0.91256025		
+	0.709	0.90730709		
+	0.7091	0.90526095		
+	0.7092	0.90199823		
+	0.7093	0.87712062		
+	0.7094	0.88347384		
+	0.7095	0.8800633		
+	0.7096	0.86066724		
+	0.7097	0.85711508		
+	0.7098	0.86923498		
+	0.7099	0.86262101		
+	0.71	0.84197031		
+	0.7101	0.84881407		
+	0.7102	0.84496974		
+	0.7103	0.85090986		
+	0.7104	0.85761862		
+	0.7105	0.86502959		
+	0.7106	0.87504876		
+	0.7107	0.88188555		
+	0.7108	0.89371229		
+	0.7109	0.90347083		
+	0.711	0.88922619		
+	0.7111	0.90267509		
+	0.7112	0.89040831		
+	0.7113	0.89565593		
+	0.7114	0.88520177		
+	0.7115	0.88247019		
+	0.7116	0.88544807		
+	0.7117	0.88708771		
+	0.7118	0.88274797		
+	0.7119	0.88034585		
+	0.712	0.86440451		
+	0.7121	0.86933393		
+	0.7122	0.866647		
+	0.7123	0.85366968		
+	0.7124	0.85649148		
+	0.7125	0.85320697		
+	0.7126	0.85901418		
+	0.7127	0.85203032		
+	0.7128	0.84859095		
+	0.7129	0.84531531		
+	0.713	0.84357551		
+	0.7131	0.84410352		
+	0.7132	0.8500366		
+	0.7133	0.8664947		
+	0.7134	0.85989097		
+	0.7135	0.86756952		
+	0.7136	0.87751447		
+	0.7137	0.8917903		
+	0.7138	0.89990655		
+	0.7139	0.89198943		
+	0.714	0.90149182		
+	0.7141	0.89640021		
+	0.7142	0.90340268		
+	0.7143	0.90008555		
+	0.7144	0.88255146		
+	0.7145	0.89392778		
+	0.7146	0.88973135		
+	0.7147	0.87294383		
+	0.7148	0.88619135		
+	0.7149	0.87909175		
+	0.715	0.87629299		
+	0.7151	0.85974398		
+	0.7152	0.87232717		
+	0.7153	0.85613547		
+	0.7154	0.85327392		
+	0.7155	0.85652828		
+	0.7156	0.86032324		
+	0.7157	0.85811631		
+	0.7158	0.84545663		
+	0.7159	0.8493264		
+	0.716	0.85644263		
+	0.7161	0.85196853		
+	0.7162	0.86148097		
+	0.7163	0.86435399		
+	0.7164	0.88676074		
+	0.7165	0.88652546		
+	0.7166	0.90135185		
+	0.7167	0.89266487		
+	0.7168	0.90020536		
+	0.7169	0.89443708		
+	0.717	0.8964443		
+	0.7171	0.90848297		
+	0.7172	0.88932885		
+	0.7173	0.89283269		
+	0.7174	0.90157838		
+	0.7175	0.90276102		
+	0.7176	0.90279822		
+	0.7177	0.89540443		
+	0.7178	0.90173212		
+	0.7179	0.89019811		
+	0.718	0.90368429		
+	0.7181	0.90187253		
+	0.7182	0.91210523		
+	0.7183	0.90722826		
+	0.7184	0.91913913		
+	0.7185	0.91646404		
+	0.7186	0.92857513		
+	0.7187	0.92150319		
+	0.7188	0.93348988		
+	0.7189	0.94199493		
+	0.719	0.93622678		
+	0.7191	0.94677039		
+	0.7192	0.9684164		
+	0.7193	0.96981992		
+	0.7194	0.98476248		
+	0.7195	1.0005337		
+	0.7196	1.0001061		
+	0.7197	1.0119511		
+	0.7198	0.99980829		
+	0.7199	1.0083149		
+	0.72	0.99650728		
+	0.7201	0.99754747		
+	0.7202	0.99119005		
+	0.7203	0.99676521		
+	0.7204	0.99967585		
+	0.7205	0.99840793		
+	0.7206	0.98736098		
+	0.7207	0.99140368		
+	0.7208	0.98197612		
+	0.7209	0.97540829		
+	0.721	0.97762417		
+	0.7211	0.97644534		
+	0.7212	0.96743603		
+	0.7213	0.96424235		
+	0.7214	0.96159416		
+	0.7215	0.96382262		
+	0.7216	0.96702275		
+	0.7217	0.95452524		
+	0.7218	0.95519849		
+	0.7219	0.96578867		
+	0.722	0.966303		
+	0.7221	0.96998225		
+	0.7222	0.99058565		
+	0.7223	1.0062906		
+	0.7224	1.002739		
+	0.7225	1.0118997		
+	0.7226	1.0251836		
+	0.7227	1.0056991		
+	0.7228	1.0152447		
+	0.7229	1.0166632		
+	0.723	1.0111905		
+	0.7231	1.0115466		
+	0.7232	0.99780204		
+	0.7233	0.99955322		
+	0.7234	0.99354774		
+	0.7235	1.0073647		
+	0.7236	0.99878993		
+	0.7237	0.9974756		
+	0.7238	0.98874876		
+	0.7239	0.974227		
+	0.724	0.9821988		
+	0.7241	0.96010602		
+	0.7242	0.97256031		
+	0.7243	0.95659119		
+	0.7244	0.95129972		
+	0.7245	0.93148769		
+	0.7246	0.93337002		
+	0.7247	0.9167904		
+	0.7248	0.91142698		
+	0.7249	0.915485		
+	0.725	0.91783316		
+	0.7251	0.92539972		
+	0.7252	0.92559472		
+	0.7253	0.93385971		
+	0.7254	0.94077625		
+	0.7255	0.92673517		
+	0.7256	0.93351874		
+	0.7257	0.92226426		
+	0.7258	0.92282459		
+	0.7259	0.91279699		
+	0.726	0.91655412		
+	0.7261	0.9120717		
+	0.7262	0.90279918		
+	0.7263	0.90546326		
+	0.7264	0.88166069		
+	0.7265	0.89373553		
+	0.7266	0.88204228		
+	0.7267	0.88152679		
+	0.7268	0.8648049		
+	0.7269	0.86390834		
+	0.727	0.85973379		
+	0.7271	0.86656652		
+	0.7272	0.84984198		
+	0.7273	0.85984691		
+	0.7274	0.84339038		
+	0.7275	0.84747912		
+	0.7276	0.84256812		
+	0.7277	0.85220697		
+	0.7278	0.85393228		
+	0.7279	0.85792204		
+	0.728	0.87281336		
+	0.7281	0.88819817		
+	0.7282	0.87973233		
+	0.7283	0.89771424		
+	0.7284	0.90257549		
+	0.7285	0.90633436		
+	0.7286	0.8973887		
+	0.7287	0.89560171		
+	0.7288	0.89721498		
+	0.7289	0.90106839		
+	0.729	0.89227742		
+	0.7291	0.88953045		
+	0.7292	0.89263263		
+	0.7293	0.8879102		
+	0.7294	0.89023791		
+	0.7295	0.87891679		
+	0.7296	0.8730626		
+	0.7297	0.86652533		
+	0.7298	0.8660776		
+	0.7299	0.86229504		
+	0.73	0.86285476		
+	0.7301	0.85764323		
+	0.7302	0.85068275		
+	0.7303	0.84559363		
+	0.7304	0.84658116		
+	0.7305	0.8457418		
+	0.7306	0.85451748		
+	0.7307	0.86424688		
+	0.7308	0.8637934		
+	0.7309	0.86008167		
+	0.731	0.87215428		
+	0.7311	0.89937846		
+	0.7312	0.90263492		
+	0.7313	0.9117421		
+	0.7314	0.90197202		
+	0.7315	0.89765824		
+	0.7316	0.91087217		
+	0.7317	0.91081089		
+	0.7318	0.89873978		
+	0.7319	0.9059204		
+	0.732	0.90574632		
+	0.7321	0.89377778		
+	0.7322	0.89761747		
+	0.7323	0.88761766		
+	0.7324	0.88659614		
+	0.7325	0.88786716		
+	0.7326	0.86587152		
+	0.7327	0.87068116		
+	0.7328	0.87285242		
+	0.7329	0.87366898		
+	0.733	0.85867279		
+	0.7331	0.85892115		
+	0.7332	0.85562906		
+	0.7333	0.84879479		
+	0.7334	0.85984981		
+	0.7335	0.85655682		
+	0.7336	0.86289384		
+	0.7337	0.86681766		
+	0.7338	0.87772139		
+	0.7339	0.88250971		
+	0.734	0.91349668		
+	0.7341	0.9245331		
+	0.7342	0.92047057		
+	0.7343	0.9366717		
+	0.7344	0.95045748		
+	0.7345	0.95399364		
+	0.7346	0.95088473		
+	0.7347	0.9498615		
+	0.7348	0.95626844		
+	0.7349	0.96367144		
+	0.735	0.95822225		
+	0.7351	0.97628411		
+	0.7352	0.96428001		
+	0.7353	0.97894235		
+	0.7354	0.97334644		
+	0.7355	0.97772473		
+	0.7356	0.97236756		
+	0.7357	0.97058102		
+	0.7358	0.97354427		
+	0.7359	0.95852199		
+	0.736	0.96475584		
+	0.7361	0.95372691		
+	0.7362	0.95377627		
+	0.7363	0.96128575		
+	0.7364	0.96728493		
+	0.7365	0.95427356		
+	0.7366	0.97267996		
+	0.7367	0.97252043		
+	0.7368	0.98271737		
+	0.7369	0.992948		
+	0.737	1.0099178		
+	0.7371	1.0164825		
+	0.7372	1.0241555		
+	0.7373	1.0121984		
+	0.7374	1.0173149		
+	0.7375	1.0148596		
+	0.7376	1.0217007		
+	0.7377	1.016574		
+	0.7378	1.0084633		
+	0.7379	1.0164296		
+	0.738	1.0070363		
+	0.7381	0.99085142		
+	0.7382	1.0003562		
+	0.7383	0.99989176		
+	0.7384	0.99822461		
+	0.7385	0.98292105		
+	0.7386	0.98816881		
+	0.7387	0.97236574		
+	0.7388	0.98396758		
+	0.7389	0.96492236		
+	0.739	0.97623156		
+	0.7391	0.96623358		
+	0.7392	0.96811351		
+	0.7393	0.96215084		
+	0.7394	0.96326888		
+	0.7395	0.96358605		
+	0.7396	0.98590506		
+	0.7397	0.98902998		
+	0.7398	0.99128234		
+	0.7399	1.0143636		
+	0.74	1.0144871		
+	0.7401	1.0205079		
+	0.7402	1.0258443		
+	0.7403	1.010268		
+	0.7404	1.0192533		
+	0.7405	0.99868027		
+	0.7406	1.0080157		
+	0.7407	0.99621943		
+	0.7408	0.98458626		
+	0.7409	0.96778765		
+	0.741	0.96826953		
+	0.7411	0.94769864		
+	0.7412	0.94135304		
+	0.7413	0.92388739		
+	0.7414	0.91426547		
+	0.7415	0.92216579		
+	0.7416	0.89702313		
+	0.7417	0.90470304		
+	0.7418	0.89068472		
+	0.7419	0.8964617		
+	0.742	0.87556699		
+	0.7421	0.87629371		
+	0.7422	0.87243717		
+	0.7423	0.86794508		
+	0.7424	0.87327674		
+	0.7425	0.87417529		
+	0.7426	0.87375823		
+	0.7427	0.89775154		
+	0.7428	0.89225387		
+	0.7429	0.91158275		
+	0.743	0.90204102		
+	0.7431	0.89912744		
+	0.7432	0.91199622		
+	0.7433	0.91168499		
+	0.7434	0.90265461		
+	0.7435	0.90326169		
+	0.7436	0.90700788		
+	0.7437	0.89990014		
+	0.7438	0.88441295		
+	0.7439	0.87878255		
+	0.744	0.89340355		
+	0.7441	0.88449936		
+	0.7442	0.88060973		
+	0.7443	0.87235058		
+	0.7444	0.87447619		
+	0.7445	0.86042622		
+	0.7446	0.87170872		
+	0.7447	0.85320257		
+	0.7448	0.85723964		
+	0.7449	0.8506655		
+	0.745	0.85337674		
+	0.7451	0.85454532		
+	0.7452	0.8527222		
+	0.7453	0.85164888		
+	0.7454	0.86073788		
+	0.7455	0.87325648		
+	0.7456	0.88552736		
+	0.7457	0.88847654		
+	0.7458	0.89042589		
+	0.7459	0.9086183		
+	0.746	0.89818607		
+	0.7461	0.91303104		
+	0.7462	0.8948492		
+	0.7463	0.89609311		
+	0.7464	0.91047517		
+	0.7465	0.90303098		
+	0.7466	0.90588454		
+	0.7467	0.89862347		
+	0.7468	0.89443616		
+	0.7469	0.88236006		
+	0.747	0.88276651		
+	0.7471	0.88527341		
+	0.7472	0.87062801		
+	0.7473	0.86327266		
+	0.7474	0.8603078		
+	0.7475	0.86063971		
+	0.7476	0.86033129		
+	0.7477	0.85237371		
+	0.7478	0.85541354		
+	0.7479	0.84881485		
+	0.748	0.85244888		
+	0.7481	0.85319465		
+	0.7482	0.85578478		
+	0.7483	0.85119793		
+	0.7484	0.86449362		
+	0.7485	0.87115351		
+	0.7486	0.89373893		
+	0.7487	0.90686347		
+	0.7488	0.89850661		
+	0.7489	0.90470233		
+	0.749	0.90397602		
+	0.7491	0.89704714		
+	0.7492	0.90774774		
+	0.7493	0.90346203		
+	0.7494	0.90327327		
+	0.7495	0.9019036		
+	0.7496	0.90652632		
+	0.7497	0.90143475		
+	0.7498	0.89660345		
+	0.7499	0.89737557		
+	0.75	0.89278976		
+	0.7501	0.88990205		
+	0.7502	0.89228933		
+	0.7503	0.88540786		
+	0.7504	0.87746868		
+	0.7505	0.88757484		
+	0.7506	0.89622357		
+	0.7507	0.89061742		
+	0.7508	0.90292573		
+	0.7509	0.90539352		
+	0.751	0.90734207		
+	0.7511	0.91345761		
+	0.7512	0.91442602		
+	0.7513	0.93107596		
+	0.7514	0.94466157		
+	0.7515	0.9699591		
+	0.7516	0.98243383		
+	0.7517	0.99187399		
+	0.7518	1.0021492		
+	0.7519	1.0009584		
+	0.752	1.0148182		
+	0.7521	1.0119195		
+	0.7522	0.99437299		
+	0.7523	0.99801069		
+	0.7524	0.99922998		
+	0.7525	1.005421		
+	0.7526	0.99078638		
+	0.7527	0.98612283		
+	0.7528	0.98878122		
+	0.7529	0.98540288		
+	0.753	0.98194179		
+	0.7531	0.97568737		
+	0.7532	0.98357161		
+	0.7533	0.98456806		
+	0.7534	0.97659599		
+	0.7535	0.9623951		
+	0.7536	0.97695206		
+	0.7537	0.95987405		
+	0.7538	0.96939389		
+	0.7539	0.97259689		
+	0.754	0.97288791		
+	0.7541	0.97229619		
+	0.7542	0.97878707		
+	0.7543	0.98379498		
+	0.7544	1.0036215		
+	0.7545	0.99997249		
+	0.7546	1.0096944		
+	0.7547	1.0180632		
+	0.7548	1.0260997		
+	0.7549	1.0251934		
+	0.755	1.0142341		
+	0.7551	1.0256548		
+	0.7552	1.0120981		
+	0.7553	1.0181692		
+	0.7554	1.0113848		
+	0.7555	1.0127836		
+	0.7556	0.9990123		
+	0.7557	1.0033256		
+	0.7558	1.0052262		
+	0.7559	0.9918986		
+	0.756	0.98173698		
+	0.7561	0.98430178		
+	0.7562	0.98511055		
+	0.7563	0.9734626		
+	0.7564	0.97873002		
+	0.7565	0.97184315		
+	0.7566	0.96380415		
+	0.7567	0.95792726		
+	0.7568	0.96077874		
+	0.7569	0.95928866		
+	0.757	0.95549591		
+	0.7571	0.9578307		
+	0.7572	0.94976959		
+	0.7573	0.94660367		
+	0.7574	0.96786434		
+	0.7575	0.96552846		
+	0.7576	0.96535753		
+	0.7577	0.94785072		
+	0.7578	0.94400645		
+	0.7579	0.94302657		
+	0.758	0.94213944		
+	0.7581	0.93098921		
+	0.7582	0.936703		
+	0.7583	0.92406725		
+	0.7584	0.91161256		
+	0.7585	0.91443079		
+	0.7586	0.90650838		
+	0.7587	0.90163218		
+	0.7588	0.88341569		
+	0.7589	0.88213165		
+	0.759	0.87776771		
+	0.7591	0.86862037		
+	0.7592	0.86633758		
+	0.7593	0.85771293		
+	0.7594	0.86589836		
+	0.7595	0.85762482		
+	0.7596	0.85352923		
+	0.7597	0.84559636		
+	0.7598	0.84297547		
+	0.7599	0.85734839		
+	0.76	0.86285227		
+	0.7601	0.85614805		
+	0.7602	0.88437689		
+	0.7603	0.88098529		
+	0.7604	0.89870147		
+	0.7605	0.91103692		
+	0.7606	0.89670152		
+	0.7607	0.90040554		
+	0.7608	0.89546703		
+	0.7609	0.89531435		
+	0.761	0.89799913		
+	0.7611	0.89814673		
+	0.7612	0.89088398		
+	0.7613	0.89695567		
+	0.7614	0.88625439		
+	0.7615	0.89395901		
+	0.7616	0.87987442		
+	0.7617	0.87928217		
+	0.7618	0.87594241		
+	0.7619	0.86623788		
+	0.762	0.87262858		
+	0.7621	0.87319537		
+	0.7622	0.85530614		
+	0.7623	0.85609013		
+	0.7624	0.8673096		
+	0.7625	0.85200304		
+	0.7626	0.84420679		
+	0.7627	0.85716363		
+	0.7628	0.85851221		
+	0.7629	0.86333225		
+	0.763	0.86089181		
+	0.7631	0.87472514		
+	0.7632	0.87491444		
+	0.7633	0.8878185		
+	0.7634	0.90493568		
+	0.7635	0.89981064		
+	0.7636	0.8986216		
+	0.7637	0.89635604		
+	0.7638	0.9111533		
+	0.7639	0.89250984		
+	0.764	0.89562748		
+	0.7641	0.89324752		
+	0.7642	0.89042833		
+	0.7643	0.88885531		
+	0.7644	0.897718		
+	0.7645	0.88235519		
+	0.7646	0.88777605		
+	0.7647	0.87725738		
+	0.7648	0.87724808		
+	0.7649	0.86967234		
+	0.765	0.86497235		
+	0.7651	0.85425951		
+	0.7652	0.86733975		
+	0.7653	0.84970295		
+	0.7654	0.85850666		
+	0.7655	0.85872824		
+	0.7656	0.85890813		
+	0.7657	0.86145508		
+	0.7658	0.85250875		
+	0.7659	0.85635834		
+	0.766	0.88154582		
+	0.7661	0.87643205		
+	0.7662	0.88631324		
+	0.7663	0.89757018		
+	0.7664	0.91037685		
+	0.7665	0.91209457		
+	0.7666	0.9109193		
+	0.7667	0.92792866		
+	0.7668	0.9222319		
+	0.7669	0.93503482		
+	0.767	0.92691567		
+	0.7671	0.93790912		
+	0.7672	0.92573834		
+	0.7673	0.94372053		
+	0.7674	0.93061875		
+	0.7675	0.93963645		
+	0.7676	0.94232915		
+	0.7677	0.94092735		
+	0.7678	0.94770183		
+	0.7679	0.95475363		
+	0.768	0.94230283		
+	0.7681	0.96138007		
+	0.7682	0.95183278		
+	0.7683	0.9480329		
+	0.7684	0.95964978		
+	0.7685	0.9636433		
+	0.7686	0.95044148		
+	0.7687	0.95877552		
+	0.7688	0.96530074		
+	0.7689	0.97780434		
+	0.769	0.98191559		
+	0.7691	0.99150899		
+	0.7692	1.0078633		
+	0.7693	1.0185791		
+	0.7694	1.0131411		
+	0.7695	1.014605		
+	0.7696	1.0134062		
+	0.7697	1.0012848		
+	0.7698	1.0076294		
+	0.7699	0.99921368		
+	0.77	1.0094051		
+	0.7701	1.0042874		
+	0.7702	0.99067875		
+	0.7703	0.99667532		
+	0.7704	0.99181229		
+	0.7705	0.98649078		
+	0.7706	0.99441175		
+	0.7707	0.98362107		
+	0.7708	0.97690265		
+	0.7709	0.97284707		
+	0.771	0.97697701		
+	0.7711	0.96587067		
+	0.7712	0.97068198		
+	0.7713	0.9763203		
+	0.7714	0.96574986		
+	0.7715	0.96725793		
+	0.7716	0.97138806		
+	0.7717	0.96687004		
+	0.7718	0.97632183		
+	0.7719	0.98010656		
+	0.772	0.9941192		
+	0.7721	1.0060866		
+	0.7722	1.0143209		
+	0.7723	1.0264518		
+	0.7724	1.0256421		
+	0.7725	1.0211827		
+	0.7726	1.024572		
+	0.7727	1.0114365		
+	0.7728	1.0064413		
+	0.7729	1.0074832		
+	0.773	1.0101438		
+	0.7731	0.99688121		
+	0.7732	0.98431826		
+	0.7733	0.9784106		
+	0.7734	0.96782081		
+	0.7735	0.95165141		
+	0.7736	0.93861694		
+	0.7737	0.93480676		
+	0.7738	0.92372044		
+	0.7739	0.92506546		
+	0.774	0.90456135		
+	0.7741	0.8978445		
+	0.7742	0.90654897		
+	0.7743	0.89030646		
+	0.7744	0.87765718		
+	0.7745	0.88391421		
+	0.7746	0.89160572		
+	0.7747	0.8927092		
+	0.7748	0.89028646		
+	0.7749	0.90298943		
+	0.775	0.91278638		
+	0.7751	0.90917181		
+	0.7752	0.91945683		
+	0.7753	0.90319105		
+	0.7754	0.91817244		
+	0.7755	0.91471937		
+	0.7756	0.89814698		
+	0.7757	0.90848909		
+	0.7758	0.90022496		
+	0.7759	0.89145471		
+	0.776	0.88878674		
+	0.7761	0.88798946		
+	0.7762	0.88034962		
+	0.7763	0.88514995		
+	0.7764	0.86373974		
+	0.7765	0.85826111		
+	0.7766	0.86127123		
+	0.7767	0.85777638		
+	0.7768	0.86011046		
+	0.7769	0.86386226		
+	0.777	0.84875871		
+	0.7771	0.84464302		
+	0.7772	0.85240538		
+	0.7773	0.84403749		
+	0.7774	0.85127887		
+	0.7775	0.85808145		
+	0.7776	0.86072115		
+	0.7777	0.87034296		
+	0.7778	0.87808568		
+	0.7779	0.88173529		
+	0.778	0.8850138		
+	0.7781	0.90173868		
+	0.7782	0.89189636		
+	0.7783	0.8960508		
+	0.7784	0.89304301		
+	0.7785	0.89355744		
+	0.7786	0.890256		
+	0.7787	0.89738441		
+	0.7788	0.8925204		
+	0.7789	0.89351306		
+	0.779	0.89215509		
+	0.7791	0.87452811		
+	0.7792	0.87346758		
+	0.7793	0.88209544		
+	0.7794	0.86218642		
+	0.7795	0.86333481		
+	0.7796	0.85798346		
+	0.7797	0.84949917		
+	0.7798	0.85310937		
+	0.7799	0.86197816		
+	0.78	0.85036414		
+	0.7801	0.84525532		
+	0.7802	0.85519123		
+	0.7803	0.84463685		
+	0.7804	0.84571205		
+	0.7805	0.86383934		
+	0.7806	0.86097173		
+	0.7807	0.88017457		
+	0.7808	0.87852033		
+	0.7809	0.8900053		
+	0.781	0.89205441		
+	0.7811	0.91065614		
+	0.7812	0.89693793		
+	0.7813	0.90663501		
+	0.7814	0.8935982		
+	0.7815	0.8865666		
+	0.7816	0.88742856		
+	0.7817	0.88326734		
+	0.7818	0.89753443		
+	0.7819	0.89075818		
+	0.782	0.88929795		
+	0.7821	0.87293702		
+	0.7822	0.8712277		
+	0.7823	0.86925144		
+	0.7824	0.87689731		
+	0.7825	0.87081662		
+	0.7826	0.86192698		
+	0.7827	0.86083737		
+	0.7828	0.86341469		
+	0.7829	0.8733669		
+	0.783	0.86887463		
+	0.7831	0.8600465		
+	0.7832	0.87417442		
+	0.7833	0.88917855		
+	0.7834	0.87979835		
+	0.7835	0.89687245		
+	0.7836	0.9218058		
+	0.7837	0.94095962		
+	0.7838	0.93844979		
+	0.7839	0.96776179		
+	0.784	0.96784897		
+	0.7841	0.9795853		
+	0.7842	0.97869255		
+	0.7843	0.97673065		
+	0.7844	0.99083186		
+	0.7845	0.9922528		
+	0.7846	0.99471915		
+	0.7847	0.99323043		
+	0.7848	0.98957089		
+	0.7849	0.97485094		
+	0.785	0.97483531		
+	0.7851	0.97754187		
+	0.7852	0.96940187		
+	0.7853	0.96552726		
+	0.7854	0.9746655		
+	0.7855	0.9650196		
+	0.7856	0.95521479		
+	0.7857	0.96607604		
+	0.7858	0.96237544		
+	0.7859	0.95855269		
+	0.786	0.96440454		
+	0.7861	0.94774096		
+	0.7862	0.95031886		
+	0.7863	0.9647559		
+	0.7864	0.96027432		
+	0.7865	0.97825894		
+	0.7866	0.98221844		
+	0.7867	1.0030759		
+	0.7868	1.0080907		
+	0.7869	1.0105879		
+	0.787	1.0039393		
+	0.7871	1.0092986		
+	0.7872	1.0055279		
+	0.7873	1.007863		
+	0.7874	0.99914403		
+	0.7875	1.0004267		
+	0.7876	1.0068571		
+	0.7877	1.0015987		
+	0.7878	0.99200846		
+	0.7879	0.98166635		
+	0.788	0.9923294		
+	0.7881	0.97303394		
+	0.7882	0.9740146		
+	0.7883	0.97053826		
+	0.7884	0.96825993		
+	0.7885	0.97043131		
+	0.7886	0.97149875		
+	0.7887	0.97254782		
+	0.7888	0.96975077		
+	0.7889	0.95252778		
+	0.789	0.96643935		
+	0.7891	0.95616532		
+	0.7892	0.95665157		
+	0.7893	0.95682541		
+	0.7894	0.96995303		
+	0.7895	0.9897334		
+	0.7896	0.98399918		
+	0.7897	0.99789933		
+	0.7898	0.98212457		
+	0.7899	0.97160606		
+	0.79	0.9756026		
+	0.7901	0.96422007		
+	0.7902	0.94971915		
+	0.7903	0.95099684		
+	0.7904	0.94525487		
+	0.7905	0.92621341		
+	0.7906	0.91952087		
+	0.7907	0.91577881		
+	0.7908	0.90432068		
+	0.7909	0.89965041		
+	0.791	0.90422487		
+	0.7911	0.88739315		
+	0.7912	0.87841429		
+	0.7913	0.87457834		
+	0.7914	0.85926701		
+	0.7915	0.85421709		
+	0.7916	0.85310304		
+	0.7917	0.85403499		
+	0.7918	0.84228898		
+	0.7919	0.85283408		
+	0.792	0.85395219		
+	0.7921	0.84293423		
+	0.7922	0.8579136		
+	0.7923	0.85641179		
+	0.7924	0.870134		
+	0.7925	0.88816049		
+	0.7926	0.89132807		
+	0.7927	0.88925343		
+	0.7928	0.89397375		
+	0.7929	0.89521665		
+	0.793	0.89010989		
+	0.7931	0.88745846		
+	0.7932	0.88249741		
+	0.7933	0.87973607		
+	0.7934	0.88516518		
+	0.7935	0.87394148		
+	0.7936	0.8815718		
+	0.7937	0.86441746		
+	0.7938	0.8728874		
+	0.7939	0.86806283		
+	0.794	0.8634056		
+	0.7941	0.85196961		
+	0.7942	0.85443318		
+	0.7943	0.85762645		
+	0.7944	0.85132678		
+	0.7945	0.85184848		
+	0.7946	0.85000663		
+	0.7947	0.85170716		
+	0.7948	0.83576208		
+	0.7949	0.83158525		
+	0.795	0.84192792		
+	0.7951	0.8559375		
+	0.7952	0.85783285		
+	0.7953	0.87504795		
+	0.7954	0.87373041		
+	0.7955	0.87814667		
+	0.7956	0.89728004		
+	0.7957	0.89485817		
+	0.7958	0.89397506		
+	0.7959	0.88708249		
+	0.796	0.88840051		
+	0.7961	0.88070157		
+	0.7962	0.89252576		
+	0.7963	0.8850929		
+	0.7964	0.87354423		
+	0.7965	0.88809476		
+	0.7966	0.87849718		
+	0.7967	0.86607987		
+	0.7968	0.8601396		
+	0.7969	0.85635922		
+	0.797	0.8615016		
+	0.7971	0.86353134		
+	0.7972	0.84495706		
+	0.7973	0.85488651		
+	0.7974	0.85493285		
+	0.7975	0.85215052		
+	0.7976	0.83916646		
+	0.7977	0.84945356		
+	0.7978	0.83204767		
+	0.7979	0.84503462		
+	0.798	0.84325751		
+	0.7981	0.84842378		
+	0.7982	0.86494503		
+	0.7983	0.88052406		
+	0.7984	0.88815834		
+	0.7985	0.88098753		
+	0.7986	0.89124214		
+	0.7987	0.90141796		
+	0.7988	0.89434412		
+	0.7989	0.90326346		
+	0.799	0.90354631		
+	0.7991	0.89593937		
+	0.7992	0.89634905		
+	0.7993	0.88704136		
+	0.7994	0.90004252		
+	0.7995	0.90293102		
+	0.7996	0.89621937		
+	0.7997	0.890949		
+	0.7998	0.9031764		
+	0.7999	0.89498996		
+	0.8	0.90973527		
+	0.8001	0.90662345		
+	0.8002	0.91588542		
+	0.8003	0.91110899		
+	0.8004	0.92430569		
+	0.8005	0.91177014		
+	0.8006	0.9172942		
+	0.8007	0.93230469		
+	0.8008	0.93877599		
+	0.8009	0.93027844		
+	0.801	0.9480144		
+	0.8011	0.95302005		
+	0.8012	0.96242017		
+	0.8013	0.9872742		
+	0.8014	0.98637577		
+	0.8015	0.99348731		
+	0.8016	0.99524688		
+	0.8017	0.98882157		
+	0.8018	0.98743763		
+	0.8019	0.9891075		
+	0.802	1.0009475		
+	0.8021	0.99922731		
+	0.8022	0.97911829		
+	0.8023	0.98249737		
+	0.8024	0.98343604		
+	0.8025	0.97556104		
+	0.8026	0.97752564		
+	0.8027	0.98205397		
+	0.8028	0.96294343		
+	0.8029	0.9700941		
+	0.803	0.95790547		
+	0.8031	0.96763596		
+	0.8032	0.95371643		
+	0.8033	0.95186602		
+	0.8034	0.9441743		
+	0.8035	0.95230742		
+	0.8036	0.94966308		
+	0.8037	0.95228926		
+	0.8038	0.94657401		
+	0.8039	0.95838944		
+	0.804	0.96735837		
+	0.8041	0.98440346		
+	0.8042	0.98534165		
+	0.8043	0.99128196		
+	0.8044	0.99108102		
+	0.8045	1.0067641		
+	0.8046	0.99310556		
+	0.8047	1.0089586		
+	0.8048	1.0090464		
+	0.8049	0.99099983		
+	0.805	0.99108733		
+	0.8051	0.9878612		
+	0.8052	0.99332143		
+	0.8053	0.99387013		
+	0.8054	0.98916105		
+	0.8055	0.98197621		
+	0.8056	0.96529271		
+	0.8057	0.97351136		
+	0.8058	0.95438997		
+	0.8059	0.95615349		
+	0.806	0.94759679		
+	0.8061	0.93887256		
+	0.8062	0.9319061		
+	0.8063	0.90994963		
+	0.8064	0.90431507		
+	0.8065	0.89472649		
+	0.8066	0.88793108		
+	0.8067	0.90016464		
+	0.8068	0.89581276		
+	0.8069	0.89823722		
+	0.807	0.89302498		
+	0.8071	0.91052515		
+	0.8072	0.91544577		
+	0.8073	0.91551772		
+	0.8074	0.90933521		
+	0.8075	0.9188098		
+	0.8076	0.9121294		
+	0.8077	0.90188281		
+	0.8078	0.88561691		
+	0.8079	0.89996814		
+	0.808	0.881292		
+	0.8081	0.88907826		
+	0.8082	0.86888457		
+	0.8083	0.87952149		
+	0.8084	0.86806576		
+	0.8085	0.85597658		
+	0.8086	0.85941173		
+	0.8087	0.86117745		
+	0.8088	0.84014727		
+	0.8089	0.84613462		
+	0.809	0.84648913		
+	0.8091	0.83059682		
+	0.8092	0.84302967		
+	0.8093	0.83077957		
+	0.8094	0.83667702		
+	0.8095	0.830074		
+	0.8096	0.83976321		
+	0.8097	0.83083781		
+	0.8098	0.84178321		
+	0.8099	0.84734223		
+	0.81	0.87269869		
+	0.8101	0.87027451		
+	0.8102	0.87648299		
+	0.8103	0.87822524		
+	0.8104	0.88214553		
+	0.8105	0.89019946		
+	0.8106	0.88763968		
+	0.8107	0.87839093		
+	0.8108	0.88375698		
+	0.8109	0.86908171		
+	0.811	0.86493077		
+	0.8111	0.86018375		
+	0.8112	0.87525934		
+	0.8113	0.85212824		
+	0.8114	0.86656178		
+	0.8115	0.84710926		
+	0.8116	0.85478817		
+	0.8117	0.83843458		
+	0.8118	0.85098011		
+	0.8119	0.83466227		
+	0.812	0.8332614		
+	0.8121	0.84408598		
+	0.8122	0.83015183		
+	0.8123	0.84015145		
+	0.8124	0.8359432		
+	0.8125	0.82501347		
+	0.8126	0.83560742		
+	0.8127	0.84241458		
+	0.8128	0.84345244		
+	0.8129	0.85577984		
+	0.813	0.8747813		
+	0.8131	0.8824426		
+	0.8132	0.87958562		
+	0.8133	0.87445925		
+	0.8134	0.87418364		
+	0.8135	0.87384161		
+	0.8136	0.8712276		
+	0.8137	0.87193191		
+	0.8138	0.88381732		
+	0.8139	0.88092121		
+	0.814	0.86422932		
+	0.8141	0.8673364		
+	0.8142	0.86800486		
+	0.8143	0.85923616		
+	0.8144	0.85598162		
+	0.8145	0.84219087		
+	0.8146	0.84045968		
+	0.8147	0.83906794		
+	0.8148	0.84045044		
+	0.8149	0.84553226		
+	0.815	0.82758583		
+	0.8151	0.84439964		
+	0.8152	0.83365535		
+	0.8153	0.8376791		
+	0.8154	0.83132988		
+	0.8155	0.83343381		
+	0.8156	0.85926453		
+	0.8157	0.87024996		
+	0.8158	0.87113198		
+	0.8159	0.88632499		
+	0.816	0.89552387		
+	0.8161	0.92187913		
+	0.8162	0.92796649		
+	0.8163	0.91773494		
+	0.8164	0.93600472		
+	0.8165	0.94319686		
+	0.8166	0.94045296		
+	0.8167	0.94257672		
+	0.8168	0.94611817		
+	0.8169	0.95404304		
+	0.817	0.94653591		
+	0.8171	0.94920838		
+	0.8172	0.9560915		
+	0.8173	0.95000098		
+	0.8174	0.93829577		
+	0.8175	0.93580902		
+	0.8176	0.94532836		
+	0.8177	0.93448872		
+	0.8178	0.93248694		
+	0.8179	0.94520281		
+	0.818	0.9289414		
+	0.8181	0.94466362		
+	0.8182	0.93129456		
+	0.8183	0.9301937		
+	0.8184	0.9462086		
+	0.8185	0.93865489		
+	0.8186	0.95041674		
+	0.8187	0.95994447		
+	0.8188	0.97780927		
+	0.8189	0.98043391		
+	0.819	0.9979261		
+	0.8191	0.99958113		
+	0.8192	0.99751311		
+	0.8193	0.99049387		
+	0.8194	0.98089114		
+	0.8195	0.99114397		
+	0.8196	0.98846879		
+	0.8197	0.98565992		
+	0.8198	0.97675318		
+	0.8199	0.98015951		
+	0.82	0.9755382		
+	0.8201	0.97457314		
+	0.8202	0.96900446		
+	0.8203	0.97001878		
+	0.8204	0.96381679		
+	0.8205	0.95467084		
+	0.8206	0.95374371		
+	0.8207	0.957918		
+	0.8208	0.95423454		
+	0.8209	0.94394864		
+	0.821	0.95136494		
+	0.8211	0.93762053		
+	0.8212	0.94939339		
+	0.8213	0.94116236		
+	0.8214	0.95006221		
+	0.8215	0.95582504		
+	0.8216	0.96688532		
+	0.8217	0.96820372		
+	0.8218	0.97795616		
+	0.8219	0.98049143		
+	0.822	0.99621679		
+	0.8221	0.99355148		
+	0.8222	0.99456678		
+	0.8223	0.98345288		
+	0.8224	0.9789395		
+	0.8225	0.96648003		
+	0.8226	0.96107407		
+	0.8227	0.94183071		
+	0.8228	0.93269842		
+	0.8229	0.92567911		
+	0.823	0.91747153		
+	0.8231	0.89517428		
+	0.8232	0.88642472		
+	0.8233	0.88972329		
+	0.8234	0.88566353		
+	0.8235	0.88072528		
+	0.8236	0.86423932		
+	0.8237	0.85871771		
+	0.8238	0.85620632		
+	0.8239	0.84676569		
+	0.824	0.83649875		
+	0.8241	0.83998867		
+	0.8242	0.83629874		
+	0.8243	0.8442493		
+	0.8244	0.85220846		
+	0.8245	0.85063478		
+	0.8246	0.8541103		
+	0.8247	0.87510469		
+	0.8248	0.8752982		
+	0.8249	0.8727875		
+	0.825	0.87845604		
+	0.8251	0.88008855		
+	0.8252	0.86967793		
+	0.8253	0.86842029		
+	0.8254	0.86222994		
+	0.8255	0.86758015		
+	0.8256	0.86579496		
+	0.8257	0.85220953		
+	0.8258	0.84648765		
+	0.8259	0.85007815		
+	0.826	0.84973161		
+	0.8261	0.84901755		
+	0.8262	0.83950641		
+	0.8263	0.84161647		
+	0.8264	0.82898495		
+	0.8265	0.83711657		
+	0.8266	0.82428878		
+	0.8267	0.82286394		
+	0.8268	0.83209297		
+	0.8269	0.82105674		
+	0.827	0.82358716		
+	0.8271	0.82033741		
+	0.8272	0.82112069		
+	0.8273	0.82822265		
+	0.8274	0.82995674		
+	0.8275	0.85375398		
+	0.8276	0.85579762		
+	0.8277	0.85939583		
+	0.8278	0.87068807		
+	0.8279	0.87326993		
+	0.828	0.87563831		
+	0.8281	0.87730098		
+	0.8282	0.87107478		
+	0.8283	0.87433507		
+	0.8284	0.86813987		
+	0.8285	0.87044693		
+	0.8286	0.85023924		
+	0.8287	0.86267477		
+	0.8288	0.85507829		
+	0.8289	0.85856619		
+	0.829	0.83774162		
+	0.8291	0.85064879		
+	0.8292	0.83611177		
+	0.8293	0.8249108		
+	0.8294	0.82304002		
+	0.8295	0.8217877		
+	0.8296	0.82281346		
+	0.8297	0.81696431		
+	0.8298	0.8324		
+	0.8299	0.82865728		
+	0.83	0.81838863		
+	0.8301	0.81373761		
+	0.8302	0.82605164		
+	0.8303	0.84353102		
+	0.8304	0.84451876		
+	0.8305	0.86259186		
+	0.8306	0.87051784		
+	0.8307	0.86533401		
+	0.8308	0.86352199		
+	0.8309	0.86774939		
+	0.831	0.86115388		
+	0.8311	0.86815587		
+	0.8312	0.87740158		
+	0.8313	0.87501254		
+	0.8314	0.86557678		
+	0.8315	0.86498135		
+	0.8316	0.85665076		
+	0.8317	0.84968152		
+	0.8318	0.85847326		
+	0.8319	0.8612971		
+	0.832	0.84813412		
+	0.8321	0.84952083		
+	0.8322	0.85914793		
+	0.8323	0.86612754		
+	0.8324	0.85977545		
+	0.8325	0.85176781		
+	0.8326	0.85495772		
+	0.8327	0.87102522		
+	0.8328	0.87217836		
+	0.8329	0.88510875		
+	0.833	0.87407308		
+	0.8331	0.8904305		
+	0.8332	0.913634		
+	0.8333	0.93102082		
+	0.8334	0.93935069		
+	0.8335	0.94814647		
+	0.8336	0.95369912		
+	0.8337	0.96062429		
+	0.8338	0.97468444		
+	0.8339	0.96939639		
+	0.834	0.96338794		
+	0.8341	0.95747382		
+	0.8342	0.96821971		
+	0.8343	0.96078045		
+	0.8344	0.97065502		
+	0.8345	0.96078382		
+	0.8346	0.9626955		
+	0.8347	0.96137569		
+	0.8348	0.95752315		
+	0.8349	0.94523575		
+	0.835	0.94775603		
+	0.8351	0.93592479		
+	0.8352	0.94393999		
+	0.8353	0.9255817		
+	0.8354	0.93974722		
+	0.8355	0.94065871		
+	0.8356	0.93227435		
+	0.8357	0.93379963		
+	0.8358	0.92870221		
+	0.8359	0.9284133		
+	0.836	0.92996965		
+	0.8361	0.94101077		
+	0.8362	0.95554516		
+	0.8363	0.95205634		
+	0.8364	0.96022752		
+	0.8365	0.97854286		
+	0.8366	0.98727722		
+	0.8367	0.97598715		
+	0.8368	0.98871198		
+	0.8369	0.96899938		
+	0.837	0.97023777		
+	0.8371	0.97673752		
+	0.8372	0.96965598		
+	0.8373	0.97879223		
+	0.8374	0.95891393		
+	0.8375	0.96720399		
+	0.8376	0.96676348		
+	0.8377	0.96221831		
+	0.8378	0.95100245		
+	0.8379	0.94017109		
+	0.838	0.94212421		
+	0.8381	0.94678106		
+	0.8382	0.92842815		
+	0.8383	0.93275634		
+	0.8384	0.9271312		
+	0.8385	0.92119344		
+	0.8386	0.92563988		
+	0.8387	0.9273609		
+	0.8388	0.9135524		
+	0.8389	0.90873838		
+	0.839	0.90658264		
+	0.8391	0.89945193		
+	0.8392	0.90468018		
+	0.8393	0.92133828		
+	0.8394	0.91416063		
+	0.8395	0.92120978		
+	0.8396	0.9093212		
+	0.8397	0.9088737		
+	0.8398	0.89603204		
+	0.8399	0.90500954		
+	0.84	0.8917844		
+	0.8401	0.88177702		
+	0.8402	0.87881147		
+	0.8403	0.8744363		
+	0.8404	0.86141448		
+	0.8405	0.86659054		
+	0.8406	0.84866527		
+	0.8407	0.85174105		
+	0.8408	0.83242663		
+	0.8409	0.84291807		
+	0.841	0.83809595		
+	0.8411	0.82200577		
+	0.8412	0.82702048		
+	0.8413	0.80966607		
+	0.8414	0.81878147		
+	0.8415	0.81858357		
+	0.8416	0.81496251		
+	0.8417	0.81643584		
+	0.8418	0.81935784		
+	0.8419	0.81515991		
+	0.842	0.82532976		
+	0.8421	0.83030929		
+	0.8422	0.84747415		
+	0.8423	0.84508293		
+	0.8424	0.85406657		
+	0.8425	0.86725385		
+	0.8426	0.86123426		
+	0.8427	0.86404914		
+	0.8428	0.85649708		
+	0.8429	0.84909222		
+	0.843	0.85548088		
+	0.8431	0.8441013		
+	0.8432	0.8429137		
+	0.8433	0.83766932		
+	0.8434	0.844795		
+	0.8435	0.8291546		
+	0.8436	0.82984451		
+	0.8437	0.83186743		
+	0.8438	0.82401075		
+	0.8439	0.82400086		
+	0.844	0.81552241		
+	0.8441	0.82697827		
+	0.8442	0.81660988		
+	0.8443	0.81042851		
+	0.8444	0.81550098		
+	0.8445	0.81351532		
+	0.8446	0.80069572		
+	0.8447	0.81801653		
+	0.8448	0.82174946		
+	0.8449	0.82584441		
+	0.845	0.82759995		
+	0.8451	0.84875123		
+	0.8452	0.85127665		
+	0.8453	0.85503467		
+	0.8454	0.85306964		
+	0.8455	0.86079177		
+	0.8456	0.86641467		
+	0.8457	0.8606129		
+	0.8458	0.86619654		
+	0.8459	0.85943433		
+	0.846	0.84859824		
+	0.8461	0.84685793		
+	0.8462	0.83706051		
+	0.8463	0.84593508		
+	0.8464	0.84681694		
+	0.8465	0.83632819		
+	0.8466	0.82594736		
+	0.8467	0.83688994		
+	0.8468	0.81847097		
+	0.8469	0.81317898		
+	0.847	0.81809924		
+	0.8471	0.82187584		
+	0.8472	0.81520213		
+	0.8473	0.80733211		
+	0.8474	0.81807203		
+	0.8475	0.81570922		
+	0.8476	0.81122946		
+	0.8477	0.80816321		
+	0.8478	0.81448674		
+	0.8479	0.82618517		
+	0.848	0.84715511		
+	0.8481	0.85134302		
+	0.8482	0.85833871		
+	0.8483	0.86235691		
+	0.8484	0.87067063		
+	0.8485	0.8750934		
+	0.8486	0.8741178		
+	0.8487	0.88508644		
+	0.8488	0.88547784		
+	0.8489	0.89346226		
+	0.849	0.89918401		
+	0.8491	0.90274475		
+	0.8492	0.89626691		
+	0.8493	0.89601049		
+	0.8494	0.89957734		
+	0.8495	0.89590146		
+	0.8496	0.90059384		
+	0.8497	0.90760706		
+	0.8498	0.91212678		
+	0.8499	0.89855428		
+	0.85	0.90889775		
+	0.8501	0.91709273		
+	0.8502	0.91369306		
+	0.8503	0.90196968		
+	0.8504	0.91053089		
+	0.8505	0.90088828		
+	0.8506	0.92029478		
+	0.8507	0.90990346		
+	0.8508	0.93159342		
+	0.8509	0.93164941		
+	0.851	0.95959667		
+	0.8511	0.9667849		
+	0.8512	0.96456614		
+	0.8513	0.97040029		
+	0.8514	0.9723414		
+	0.8515	0.9729969		
+	0.8516	0.95705686		
+	0.8517	0.95629695		
+	0.8518	0.96796878		
+	0.8519	0.96074107		
+	0.852	0.96337323		
+	0.8521	0.949379		
+	0.8522	0.93927719		
+	0.8523	0.9403256		
+	0.8524	0.93178366		
+	0.8525	0.94418835		
+	0.8526	0.92653781		
+	0.8527	0.92409666		
+	0.8528	0.93067637		
+	0.8529	0.92104442		
+	0.853	0.93105105		
+	0.8531	0.92606537		
+	0.8532	0.9271276		
+	0.8533	0.92587354		
+	0.8534	0.91767822		
+	0.8535	0.91864379		
+	0.8536	0.92312599		
+	0.8537	0.9416233		
+	0.8538	0.94192117		
+	0.8539	0.96348591		
+	0.854	0.95382883		
+	0.8541	0.95978906		
+	0.8542	0.97387529		
+	0.8543	0.97985973		
+	0.8544	0.95981126		
+	0.8545	0.95843388		
+	0.8546	0.95431977		
+	0.8547	0.97040517		
+	0.8548	0.94860692		
+	0.8549	0.95851231		
+	0.855	0.95448825		
+	0.8551	0.9408863		
+	0.8552	0.93108523		
+	0.8553	0.91432867		
+	0.8554	0.91403933		
+	0.8555	0.89999946		
+	0.8556	0.88469715		
+	0.8557	0.87062857		
+	0.8558	0.86740339		
+	0.8559	0.85612775		
+	0.856	0.85564604		
+	0.8561	0.83750287		
+	0.8562	0.8425419		
+	0.8563	0.83845885		
+	0.8564	0.82479567		
+	0.8565	0.83465635		
+	0.8566	0.83745943		
+	0.8567	0.8441155		
+	0.8568	0.84510164		
+	0.8569	0.85172087		
+	0.857	0.86034469		
+	0.8571	0.86936947		
+	0.8572	0.85305192		
+	0.8573	0.85791531		
+	0.8574	0.86439721		
+	0.8575	0.86180672		
+	0.8576	0.84447909		
+	0.8577	0.84782568		
+	0.8578	0.84484954		
+	0.8579	0.82991209		
+	0.858	0.84320231		
+	0.8581	0.83686329		
+	0.8582	0.82844505		
+	0.8583	0.81754628		
+	0.8584	0.81969019		
+	0.8585	0.81863468		
+	0.8586	0.80411297		
+	0.8587	0.81171938		
+	0.8588	0.80408731		
+	0.8589	0.81045579		
+	0.859	0.80294453		
+	0.8591	0.79860795		
+	0.8592	0.79322711		
+	0.8593	0.80205003		
+	0.8594	0.80188848		
+	0.8595	0.80127873		
+	0.8596	0.82015959		
+	0.8597	0.8263385		
+	0.8598	0.84700454		
+	0.8599	0.84925785		
+	0.86	0.84911791		
+	0.8601	0.86074844		
+	0.8602	0.85094968		
+	0.8603	0.84416475		
+	0.8604	0.84387669		
+	0.8605	0.84373751		
+	0.8606	0.8475806		
+	0.8607	0.84748077		
+	0.8608	0.83972109		
+	0.8609	0.83368527		
+	0.861	0.82346743		
+	0.8611	0.82178351		
+	0.8612	0.81797908		
+	0.8613	0.81688987		
+	0.8614	0.81229214		
+	0.8615	0.81646104		
+	0.8616	0.79802474		
+	0.8617	0.80028799		
+	0.8618	0.81060243		
+	0.8619	0.80540878		
+	0.862	0.80130666		
+	0.8621	0.80394992		
+	0.8622	0.79913717		
+	0.8623	0.796549		
+	0.8624	0.80520279		
+	0.8625	0.81309172		
+	0.8626	0.83680615		
+	0.8627	0.83117064		
+	0.8628	0.84116945		
+	0.8629	0.84917116		
+	0.863	0.85699139		
+	0.8631	0.85455736		
+	0.8632	0.85797773		
+	0.8633	0.84260967		
+	0.8634	0.83637495		
+	0.8635	0.83639002		
+	0.8636	0.83805564		
+	0.8637	0.82849475		
+	0.8638	0.84165467		
+	0.8639	0.84030186		
+	0.864	0.83385403		
+	0.8641	0.83005755		
+	0.8642	0.82006519		
+	0.8643	0.82411214		
+	0.8644	0.81516295		
+	0.8645	0.81202126		
+	0.8646	0.8208701		
+	0.8647	0.8134268		
+	0.8648	0.8183695		
+	0.8649	0.81132432		
+	0.865	0.82271136		
+	0.8651	0.82825914		
+	0.8652	0.82911146		
+	0.8653	0.84829782		
+	0.8654	0.85849743		
+	0.8655	0.8726018		
+	0.8656	0.88996899		
+	0.8657	0.90270903		
+	0.8658	0.91995762		
+	0.8659	0.92226328		
+	0.866	0.92891187		
+	0.8661	0.92588592		
+	0.8662	0.92956917		
+	0.8663	0.94547317		
+	0.8664	0.92949103		
+	0.8665	0.9454401		
+	0.8666	0.93767733		
+	0.8667	0.9313519		
+	0.8668	0.93051617		
+	0.8669	0.92506088		
+	0.867	0.91484983		
+	0.8671	0.92567065		
+	0.8672	0.91728565		
+	0.8673	0.90871215		
+	0.8674	0.92111633		
+	0.8675	0.91560835		
+	0.8676	0.90525823		
+	0.8677	0.9055144		
+	0.8678	0.911668		
+	0.8679	0.91038247		
+	0.868	0.9001275		
+	0.8681	0.90886114		
+	0.8682	0.91737613		
+	0.8683	0.92118999		
+	0.8684	0.92883607		
+	0.8685	0.95118432		
+	0.8686	0.94751654		
+	0.8687	0.94809563		
+	0.8688	0.9607321		
+	0.8689	0.96870253		
+	0.869	0.96141681		
+	0.8691	0.96651404		
+	0.8692	0.96485676		
+	0.8693	0.95640004		
+	0.8694	0.96106084		
+	0.8695	0.94896822		
+	0.8696	0.94838365		
+	0.8697	0.93979421		
+	0.8698	0.94457764		
+	0.8699	0.94060414		
+	0.87	0.92875297		
+	0.8701	0.9340941		
+	0.8702	0.92170455		
+	0.8703	0.91734164		
+	0.8704	0.92059515		
+	0.8705	0.91775533		
+	0.8706	0.90594493		
+	0.8707	0.91257755		
+	0.8708	0.9031878		
+	0.8709	0.90509233		
+	0.871	0.89812753		
+	0.8711	0.90779892		
+	0.8712	0.92084144		
+	0.8713	0.93340561		
+	0.8714	0.93107805		
+	0.8715	0.92876608		
+	0.8716	0.94022263		
+	0.8717	0.93868013		
+	0.8718	0.92914246		
+	0.8719	0.92696355		
+	0.872	0.90413435		
+	0.8721	0.90162613		
+	0.8722	0.9016331		
+	0.8723	0.88546784		
+	0.8724	0.89098286		
+	0.8725	0.87692575		
+	0.8726	0.86491781		
+	0.8727	0.86133428		
+	0.8728	0.85160999		
+	0.8729	0.84576892		
+	0.873	0.84353803		
+	0.8731	0.83479162		
+	0.8732	0.8194119		
+	0.8733	0.81445192		
+	0.8734	0.80714667		
+	0.8735	0.81573437		
+	0.8736	0.80551428		
+	0.8737	0.79291149		
+	0.8738	0.79692723		
+	0.8739	0.7872245		
+	0.874	0.78950017		
+	0.8741	0.79941734		
+	0.8742	0.81769513		
+	0.8743	0.81223269		
+	0.8744	0.83614263		
+	0.8745	0.83442627		
+	0.8746	0.84999857		
+	0.8747	0.83753499		
+	0.8748	0.84403155		
+	0.8749	0.8302163		
+	0.875	0.84343836		
+	0.8751	0.82779523		
+	0.8752	0.84010431		
+	0.8753	0.83768943		
+	0.8754	0.83416327		
+	0.8755	0.82699429		
+	0.8756	0.82428608		
+	0.8757	0.80738131		
+	0.8758	0.82304203		
+	0.8759	0.81754862		
+	0.876	0.81005032		
+	0.8761	0.81154869		
+	0.8762	0.79286753		
+	0.8763	0.8047235		
+	0.8764	0.79365569		
+	0.8765	0.79365981		
+	0.8766	0.79773425		
+	0.8767	0.78457891		
+	0.8768	0.79269053		
+	0.8769	0.79776701		
+	0.877	0.79402921		
+	0.8771	0.8003969		
+	0.8772	0.81390348		
+	0.8773	0.82635626		
+	0.8774	0.82843649		
+	0.8775	0.83915278		
+	0.8776	0.83648959		
+	0.8777	0.8390246		
+	0.8778	0.83180238		
+	0.8779	0.83030115		
+	0.878	0.84110648		
+	0.8781	0.83625393		
+	0.8782	0.82623478		
+	0.8783	0.82442084		
+	0.8784	0.82780885		
+	0.8785	0.82199028		
+	0.8786	0.81170481		
+	0.8787	0.80746575		
+	0.8788	0.81790129		
+	0.8789	0.8041376		
+	0.879	0.80695636		
+	0.8791	0.7954182		
+	0.8792	0.80051809		
+	0.8793	0.78798631		
+	0.8794	0.78632408		
+	0.8795	0.79694139		
+	0.8796	0.79367674		
+	0.8797	0.79590766		
+	0.8798	0.78844651		
+	0.8799	0.79595071		
+	0.88	0.80522878		
+	0.8801	0.81440379		
+	0.8802	0.82378646		
+	0.8803	0.82639758		
+	0.8804	0.8484825		
+	0.8805	0.83933957		
+	0.8806	0.84563882		
+	0.8807	0.84372068		
+	0.8808	0.8532521		
+	0.8809	0.85370699		
+	0.881	0.85474176		
+	0.8811	0.83674491		
+	0.8812	0.85530103		
+	0.8813	0.85367755		
+	0.8814	0.84869782		
+	0.8815	0.85441751		
+	0.8816	0.85838082		
+	0.8817	0.85900883		
+	0.8818	0.85963853		
+	0.8819	0.84662329		
+	0.882	0.86393064		
+	0.8821	0.86008739		
+	0.8822	0.86720959		
+	0.8823	0.87576427		
+	0.8824	0.86455666		
+	0.8825	0.87561455		
+	0.8826	0.87085595		
+	0.8827	0.87610354		
+	0.8828	0.879102		
+	0.8829	0.90774751		
+	0.883	0.90198003		
+	0.8831	0.92934238		
+	0.8832	0.92206786		
+	0.8833	0.93923763		
+	0.8834	0.95010751		
+	0.8835	0.94099868		
+	0.8836	0.9441344		
+	0.8837	0.9419714		
+	0.8838	0.93930236		
+	0.8839	0.94621424		
+	0.884	0.94381636		
+	0.8841	0.94313603		
+	0.8842	0.94026422		
+	0.8843	0.9225461		
+	0.8844	0.92090127		
+	0.8845	0.92798599		
+	0.8846	0.92679101		
+	0.8847	0.90789381		
+	0.8848	0.91532893		
+	0.8849	0.91976981		
+	0.885	0.90645381		
+	0.8851	0.90592055		
+	0.8852	0.89569545		
+	0.8853	0.91270738		
+	0.8854	0.89777358		
+	0.8855	0.90919705		
+	0.8856	0.90902387		
+	0.8857	0.89858318		
+	0.8858	0.91188556		
+	0.8859	0.92717627		
+	0.886	0.92466291		
+	0.8861	0.93039288		
+	0.8862	0.9374191		
+	0.8863	0.95894941		
+	0.8864	0.94304732		
+	0.8865	0.94999252		
+	0.8866	0.94588226		
+	0.8867	0.94410989		
+	0.8868	0.95056877		
+	0.8869	0.93645651		
+	0.887	0.93636052		
+	0.8871	0.94629652		
+	0.8872	0.93546464		
+	0.8873	0.92458466		
+	0.8874	0.93418002		
+	0.8875	0.92339215		
+	0.8876	0.92592847		
+	0.8877	0.91238052		
+	0.8878	0.89572331		
+	0.8879	0.89195205		
+	0.888	0.89369541		
+	0.8881	0.88301142		
+	0.8882	0.86020168		
+	0.8883	0.85858094		
+	0.8884	0.84789134		
+	0.8885	0.84824389		
+	0.8886	0.83448336		
+	0.8887	0.84541058		
+	0.8888	0.85162823		
+	0.8889	0.85467562		
+	0.889	0.85972315		
+	0.8891	0.86697545		
+	0.8892	0.87184311		
+	0.8893	0.86602752		
+	0.8894	0.86470905		
+	0.8895	0.86230319		
+	0.8896	0.85695085		
+	0.8897	0.83975769		
+	0.8898	0.83978327		
+	0.8899	0.8450677		
+	0.89	0.83554073		
+	0.8901	0.83560618		
+	0.8902	0.81429115		
+	0.8903	0.82188875		
+	0.8904	0.8114818		
+	0.8905	0.81300293		
+	0.8906	0.79259329		
+	0.8907	0.80058079		
+	0.8908	0.78525574		
+	0.8909	0.79861233		
+	0.891	0.79848726		
+	0.8911	0.79487704		
+	0.8912	0.79080931		
+	0.8913	0.774921		
+	0.8914	0.78754512		
+	0.8915	0.77958706		
+	0.8916	0.78555683		
+	0.8917	0.8028638		
+	0.8918	0.80613204		
+	0.8919	0.81719395		
+	0.892	0.81807162		
+	0.8921	0.82577351		
+	0.8922	0.83118965		
+	0.8923	0.83392315		
+	0.8924	0.83997687		
+	0.8925	0.8300416		
+	0.8926	0.83939611		
+	0.8927	0.8201334		
+	0.8928	0.82290596		
+	0.8929	0.82483871		
+	0.893	0.82415104		
+	0.8931	0.82456174		
+	0.8932	0.80387025		
+	0.8933	0.81682618		
+	0.8934	0.79913767		
+	0.8935	0.79424179		
+	0.8936	0.80180694		
+	0.8937	0.79317214		
+	0.8938	0.79845903		
+	0.8939	0.78361839		
+	0.894	0.78043456		
+	0.8941	0.79498952		
+	0.8942	0.78120145		
+	0.8943	0.78104087		
+	0.8944	0.78981009		
+	0.8945	0.79254886		
+	0.8946	0.79340674		
+	0.8947	0.80759607		
+	0.8948	0.81107627		
+	0.8949	0.81727799		
+	0.895	0.83688919		
+	0.8951	0.84514957		
+	0.8952	0.83526773		
+	0.8953	0.83585784		
+	0.8954	0.82943833		
+	0.8955	0.8335478		
+	0.8956	0.82666132		
+	0.8957	0.8365008		
+	0.8958	0.82363859		
+	0.8959	0.82148738		
+	0.896	0.82023711		
+	0.8961	0.81931343		
+	0.8962	0.80595895		
+	0.8963	0.8001243		
+	0.8964	0.79463746		
+	0.8965	0.80730414		
+	0.8966	0.80027203		
+	0.8967	0.795943		
+	0.8968	0.79062876		
+	0.8969	0.79421584		
+	0.897	0.78496873		
+	0.8971	0.79742528		
+	0.8972	0.79042372		
+	0.8973	0.78695464		
+	0.8974	0.79688196		
+	0.8975	0.80577987		
+	0.8976	0.81778054		
+	0.8977	0.83527009		
+	0.8978	0.84127631		
+	0.8979	0.86173271		
+	0.898	0.8648261		
+	0.8981	0.88389241		
+	0.8982	0.87540264		
+	0.8983	0.87603748		
+	0.8984	0.88308182		
+	0.8985	0.89719968		
+	0.8986	0.89879625		
+	0.8987	0.89462386		
+	0.8988	0.89102805		
+	0.8989	0.90488029		
+	0.899	0.90142595		
+	0.8991	0.8967472		
+	0.8992	0.90756112		
+	0.8993	0.90098264		
+	0.8994	0.89014747		
+	0.8995	0.89278119		
+	0.8996	0.89907723		
+	0.8997	0.89763188		
+	0.8998	0.90039467		
+	0.8999	0.88216694		
+	0.9	0.88329718		
+	0.9001	0.89398437		
+	0.9002	0.89693485		
+	0.9003	0.8851608		
+	0.9004	0.89533869		
+	0.9005	0.90887386		
+	0.9006	0.91580535		
+	0.9007	0.92844252		
+	0.9008	0.93684965		
+	0.9009	0.94874035		
+	0.901	0.94072585		
+	0.9011	0.93856521		
+	0.9012	0.94263215		
+	0.9013	0.94423131		
+	0.9014	0.94439377		
+	0.9015	0.93043999		
+	0.9016	0.9375783		
+	0.9017	0.93903335		
+	0.9018	0.935459		
+	0.9019	0.92454855		
+	0.902	0.92273965		
+	0.9021	0.91160559		
+	0.9022	0.91622443		
+	0.9023	0.90938986		
+	0.9024	0.90435564		
+	0.9025	0.90896849		
+	0.9026	0.89257985		
+	0.9027	0.90482172		
+	0.9028	0.90540228		
+	0.9029	0.89274264		
+	0.903	0.88629836		
+	0.9031	0.9026903		
+	0.9032	0.90107673		
+	0.9033	0.89963798		
+	0.9034	0.92088772		
+	0.9035	0.92245381		
+	0.9036	0.93466635		
+	0.9037	0.93173343		
+	0.9038	0.9462505		
+	0.9039	0.93717225		
+	0.904	0.95417447		
+	0.9041	0.93641995		
+	0.9042	0.93381917		
+	0.9043	0.93250888		
+	0.9044	0.92721161		
+	0.9045	0.90545638		
+	0.9046	0.90281829		
+	0.9047	0.88856409		
+	0.9048	0.88980861		
+	0.9049	0.87747216		
+	0.905	0.86807029		
+	0.9051	0.85664511		
+	0.9052	0.83652477		
+	0.9053	0.8330466		
+	0.9054	0.83024728		
+	0.9055	0.81843989		
+	0.9056	0.82184251		
+	0.9057	0.80950853		
+	0.9058	0.80829073		
+	0.9059	0.79208514		
+	0.906	0.79515002		
+	0.9061	0.79595289		
+	0.9062	0.79263709		
+	0.9063	0.81269526		
+	0.9064	0.80823059		
+	0.9065	0.82211838		
+	0.9066	0.82262454		
+	0.9067	0.82418357		
+	0.9068	0.83638791		
+	0.9069	0.8386135		
+	0.907	0.83516236		
+	0.9071	0.836536		
+	0.9072	0.83161806		
+	0.9073	0.83514035		
+	0.9074	0.81741933		
+	0.9075	0.81536125		
+	0.9076	0.81387021		
+	0.9077	0.8109914		
+	0.9078	0.80256466		
+	0.9079	0.80091987		
+	0.908	0.79640524		
+	0.9081	0.79649521		
+	0.9082	0.7934718		
+	0.9083	0.78735505		
+	0.9084	0.79250852		
+	0.9085	0.77978181		
+	0.9086	0.79250741		
+	0.9087	0.7822321		
+	0.9088	0.79026016		
+	0.9089	0.77158346		
+	0.909	0.78811016		
+	0.9091	0.7799595		
+	0.9092	0.79216311		
+	0.9093	0.79430139		
+	0.9094	0.82079382		
+	0.9095	0.81796997		
+	0.9096	0.83507404		
+	0.9097	0.8320921		
+	0.9098	0.83430241		
+	0.9099	0.82766533		
+	0.91	0.83984205		
+	0.9101	0.82012495		
+	0.9102	0.82332784		
+	0.9103	0.82883449		
+	0.9104	0.81831538		
+	0.9105	0.8186996		
+	0.9106	0.80664905		
+	0.9107	0.81450602		
+	0.9108	0.79908538		
+	0.9109	0.80534121		
+	0.911	0.79552302		
+	0.9111	0.80390426		
+	0.9112	0.79929002		
+	0.9113	0.7906346		
+	0.9114	0.79108976		
+	0.9115	0.78876169		
+	0.9116	0.79217742		
+	0.9117	0.77673982		
+	0.9118	0.79037325		
+	0.9119	0.77963123		
+	0.912	0.78480829		
+	0.9121	0.78227113		
+	0.9122	0.79678125		
+	0.9123	0.80984666		
+	0.9124	0.8164841		
+	0.9125	0.82541617		
+	0.9126	0.83444619		
+	0.9127	0.83700277		
+	0.9128	0.84091503		
+	0.9129	0.82456086		
+	0.913	0.82965299		
+	0.9131	0.83318041		
+	0.9132	0.82073751		
+	0.9133	0.81803267		
+	0.9134	0.82139846		
+	0.9135	0.82589481		
+	0.9136	0.82655837		
+	0.9137	0.82711509		
+	0.9138	0.80929057		
+	0.9139	0.81082389		
+	0.914	0.81827469		
+	0.9141	0.80648321		
+	0.9142	0.80898703		
+	0.9143	0.82772323		
+	0.9144	0.8299866		
+	0.9145	0.83108982		
+	0.9146	0.8242618		
+	0.9147	0.83936761		
+	0.9148	0.82942693		
+	0.9149	0.84462933		
+	0.915	0.86368593		
+	0.9151	0.86991464		
+	0.9152	0.89466751		
+	0.9153	0.90024517		
+	0.9154	0.90891273		
+	0.9155	0.92446014		
+	0.9156	0.93026761		
+	0.9157	0.92907817		
+	0.9158	0.92494376		
+	0.9159	0.93344988		
+	0.916	0.93779652		
+	0.9161	0.9290801		
+	0.9162	0.92872263		
+	0.9163	0.92091337		
+	0.9164	0.91892567		
+	0.9165	0.911519		
+	0.9166	0.91611391		
+	0.9167	0.90650661		
+	0.9168	0.91415726		
+	0.9169	0.90816312		
+	0.917	0.89877113		
+	0.9171	0.90335002		
+	0.9172	0.89133482		
+	0.9173	0.90530965		
+	0.9174	0.89026419		
+	0.9175	0.89690063		
+	0.9176	0.8901009		
+	0.9177	0.88258384		
+	0.9178	0.90363273		
+	0.9179	0.90185024		
+	0.918	0.91353139		
+	0.9181	0.91457803		
+	0.9182	0.92559301		
+	0.9183	0.94072963		
+	0.9184	0.94762642		
+	0.9185	0.94376858		
+	0.9186	0.95405884		
+	0.9187	0.94857919		
+	0.9188	0.94645487		
+	0.9189	0.94673979		
+	0.919	0.9488685		
+	0.9191	0.93885031		
+	0.9192	0.92912489		
+	0.9193	0.93839499		
+	0.9194	0.92635369		
+	0.9195	0.92295251		
+	0.9196	0.9124146		
+	0.9197	0.91250535		
+	0.9198	0.91371726		
+	0.9199	0.91124576		
+	0.92	0.90060247		
+	0.9201	0.90782848		
+	0.9202	0.90211768		
+	0.9203	0.89526528		
+	0.9204	0.88744372		
+	0.9205	0.88480413		
+	0.9206	0.88999421		
+	0.9207	0.88593049		
+	0.9208	0.87870546		
+	0.9209	0.88519298		
+	0.921	0.87453643		
+	0.9211	0.87997165		
+	0.9212	0.88197556		
+	0.9213	0.89804172		
+	0.9214	0.89475703		
+	0.9215	0.87954725		
+	0.9216	0.88240709		
+	0.9217	0.86993808		
+	0.9218	0.8725663		
+	0.9219	0.86656002		
+	0.922	0.85411194		
+	0.9221	0.85392367		
+	0.9222	0.83638568		
+	0.9223	0.83501567		
+	0.9224	0.83249111		
+	0.9225	0.82471516		
+	0.9226	0.82441787		
+	0.9227	0.80683901		
+	0.9228	0.81114443		
+	0.9229	0.80800135		
+	0.923	0.80021811		
+	0.9231	0.79903902		
+	0.9232	0.79075689		
+	0.9233	0.78911334		
+	0.9234	0.77393415		
+	0.9235	0.7838775		
+	0.9236	0.78651103		
+	0.9237	0.77391176		
+	0.9238	0.78540285		
+	0.9239	0.8056472		
+	0.924	0.81429839		
+	0.9241	0.81075242		
+	0.9242	0.81923745		
+	0.9243	0.83509013		
+	0.9244	0.83468165		
+	0.9245	0.83963122		
+	0.9246	0.83922347		
+	0.9247	0.82329035		
+	0.9248	0.82391599		
+	0.9249	0.81673887		
+	0.925	0.81944103		
+	0.9251	0.81614162		
+	0.9252	0.81071671		
+	0.9253	0.82012759		
+	0.9254	0.80560817		
+	0.9255	0.81050582		
+	0.9256	0.79495439		
+	0.9257	0.78869915		
+	0.9258	0.7959944		
+	0.9259	0.79697349		
+	0.926	0.77909746		
+	0.9261	0.7777416		
+	0.9262	0.78864794		
+	0.9263	0.79114711		
+	0.9264	0.78273927		
+	0.9265	0.77247273		
+	0.9266	0.7750521		
+	0.9267	0.79176488		
+	0.9268	0.80419273		
+	0.9269	0.80431663		
+	0.927	0.81134574		
+	0.9271	0.83463761		
+	0.9272	0.83314879		
+	0.9273	0.84282212		
+	0.9274	0.83768972		
+	0.9275	0.82800447		
+	0.9276	0.8244628		
+	0.9277	0.83141569		
+	0.9278	0.82063407		
+	0.9279	0.82919375		
+	0.928	0.81858572		
+	0.9281	0.80890769		
+	0.9282	0.8169637		
+	0.9283	0.80710955		
+	0.9284	0.80095054		
+	0.9285	0.8121643		
+	0.9286	0.80059201		
+	0.9287	0.78967913		
+	0.9288	0.79000298		
+	0.9289	0.79609767		
+	0.929	0.78160857		
+	0.9291	0.78696277		
+	0.9292	0.78254748		
+	0.9293	0.77480419		
+	0.9294	0.78089372		
+	0.9295	0.77955287		
+	0.9296	0.79829918		
+	0.9297	0.7936081		
+	0.9298	0.81165018		
+	0.9299	0.81840026		
+	0.93	0.83860428		
+	0.9301	0.84424801		
+	0.9302	0.83783625		
+	0.9303	0.85352923		
+	0.9304	0.85771689		
+	0.9305	0.85136725		
+	0.9306	0.86316997		
+	0.9307	0.86602201		
+	0.9308	0.85785029		
+	0.9309	0.85567315		
+	0.931	0.8614579		
+	0.9311	0.8754589		
+	0.9312	0.86914531		
+	0.9313	0.87024622		
+	0.9314	0.87811903		
+	0.9315	0.86603656		
+	0.9316	0.87128445		
+	0.9317	0.88445411		
+	0.9318	0.88888014		
+	0.9319	0.87131676		
+	0.932	0.88239995		
+	0.9321	0.87628878		
+	0.9322	0.87468598		
+	0.9323	0.8738901		
+	0.9324	0.88181556		
+	0.9325	0.88910211		
+	0.9326	0.89676197		
+	0.9327	0.90233095		
+	0.9328	0.92650437		
+	0.9329	0.93174826		
+	0.933	0.92966577		
+	0.9331	0.92998293		
+	0.9332	0.94317712		
+	0.9333	0.93638325		
+	0.9334	0.9311788		
+	0.9335	0.93088317		
+	0.9336	0.94524365		
+	0.9337	0.92984305		
+	0.9338	0.93006843		
+	0.9339	0.92810884		
+	0.934	0.92589308		
+	0.9341	0.9234937		
+	0.9342	0.92219135		
+	0.9343	0.92506609		
+	0.9344	0.91937065		
+	0.9345	0.90650719		
+	0.9346	0.90727129		
+	0.9347	0.89631926		
+	0.9348	0.89958787		
+	0.9349	0.90220234		
+	0.935	0.89839564		
+	0.9351	0.89773967		
+	0.9352	0.88694892		
+	0.9353	0.90463921		
+	0.9354	0.88975065		
+	0.9355	0.89723507		
+	0.9356	0.91727961		
+	0.9357	0.92995069		
+	0.9358	0.92694798		
+	0.9359	0.94947455		
+	0.936	0.94759176		
+	0.9361	0.94617676		
+	0.9362	0.95427938		
+	0.9363	0.94359849		
+	0.9364	0.93778143		
+	0.9365	0.94456955		
+	0.9366	0.93911531		
+	0.9367	0.93061345		
+	0.9368	0.92896076		
+	0.9369	0.92357001		
+	0.937	0.91953756		
+	0.9371	0.91054679		
+	0.9372	0.91257673		
+	0.9373	0.89459343		
+	0.9374	0.87500756		
+	0.9375	0.87840881		
+	0.9376	0.85330034		
+	0.9377	0.85387099		
+	0.9378	0.84578743		
+	0.9379	0.83036574		
+	0.938	0.82929222		
+	0.9381	0.8186571		
+	0.9382	0.82275171		
+	0.9383	0.82384175		
+	0.9384	0.83129552		
+	0.9385	0.82505832		
+	0.9386	0.8432904		
+	0.9387	0.84380571		
+	0.9388	0.84465629		
+	0.9389	0.8515928		
+	0.939	0.84215317		
+	0.9391	0.85264525		
+	0.9392	0.83247305		
+	0.9393	0.84609468		
+	0.9394	0.8348202		
+	0.9395	0.8330395		
+	0.9396	0.82919346		
+	0.9397	0.83237329		
+	0.9398	0.81233441		
+	0.9399	0.81579882		
+	0.94	0.81021276		
+	0.9401	0.80273006		
+	0.9402	0.80261588		
+	0.9403	0.80649984		
+	0.9404	0.79930496		
+	0.9405	0.79040666		
+	0.9406	0.79993319		
+	0.9407	0.78783291		
+	0.9408	0.79463473		
+	0.9409	0.79050312		
+	0.941	0.77549401		
+	0.9411	0.77342738		
+	0.9412	0.78926269		
+	0.9413	0.79446115		
+	0.9414	0.79218834		
+	0.9415	0.80907722		
+	0.9416	0.81813526		
+	0.9417	0.82253708		
+	0.9418	0.84156752		
+	0.9419	0.83944712		
+	0.942	0.84548094		
+	0.9421	0.84419418		
+	0.9422	0.84277083		
+	0.9423	0.83061214		
+	0.9424	0.82471389		
+	0.9425	0.82136099		
+	0.9426	0.8286088		
+	0.9427	0.81396653		
+	0.9428	0.81249319		
+	0.9429	0.82061765		
+	0.943	0.81158959		
+	0.9431	0.81020215		
+	0.9432	0.80373809		
+	0.9433	0.80199159		
+	0.9434	0.79144172		
+	0.9435	0.79181161		
+	0.9436	0.79868922		
+	0.9437	0.78333889		
+	0.9438	0.78103792		
+	0.9439	0.78102099		
+	0.944	0.78756841		
+	0.9441	0.78809119		
+	0.9442	0.78336531		
+	0.9443	0.79377079		
+	0.9444	0.80817537		
+	0.9445	0.8114884		
+	0.9446	0.82571633		
+	0.9447	0.84160515		
+	0.9448	0.83681112		
+	0.9449	0.83138448		
+	0.945	0.83813547		
+	0.9451	0.8377067		
+	0.9452	0.8434897		
+	0.9453	0.82496732		
+	0.9454	0.82242445		
+	0.9455	0.8348596		
+	0.9456	0.82409857		
+	0.9457	0.81384489		
+	0.9458	0.80956924		
+	0.9459	0.81968419		
+	0.946	0.8131374		
+       r       0				
.ends				
