.subckt ori n1 n2				
vin n1 n2 pwl				
+	0.0001	0.207		
+	0.0002	0.81		
+	0.0003	1.805		
+	0.0004	3.267		
+	0.0005	5.32		
+	0.0006	8.026		
+	0.0007	11.385		
+	0.0008	15.129		
+	0.0009	19.123		
+	0.001	23.508		
+	0.0011	28.534		
+	0.0012	33.622		
+	0.0013	39.071		
+	0.0014	45.211		
+	0.0015	51.493		
+	0.0016	57.943		
+	0.0017	64.661		
+	0.0018	71.448		
+	0.0019	77.998		
+	0.002	84.286		
+	0.0021	89.773		
+	0.0022	93.803		
+	0.0023	96.739		
+	0.0024	99.004		
+	0.0025	100.49		
+	0.0026	101.38		
+	0.0027	102.039		
+	0.0028	102.593		
+	0.0029	102.922		
+	0.003	103.482		
+	0.0031	104.135		
+	0.0032	104.745		
+	0.0033	105.473		
+	0.0034	106.381		
+	0.0035	107.245		
+	0.0036	107.874		
+	0.0037	108.72		
+	0.0038	109.366		
+	0.0039	109.796		
+	0.004	110.237		
+	0.0041	110.685		
+	0.0042	111.009		
+	0.0043	111.096		
+	0.0044	111.345		
+	0.0045	111.519		
+	0.0046	111.5		
+	0.0047	111.631		
+	0.0048	111.824		
+	0.0049	111.656		
+	0.005	111.724		
+	0.0051	111.805		
+	0.0052	111.792		
+	0.0053	111.736		
+	0.0054	111.83		
+	0.0055	111.836		
+	0.0056	111.699		
+	0.0057	111.749		
+	0.0058	111.979		
+	0.0059	111.898		
+	0.006	112.004		
+	0.0061	112.315		
+	0.0062	112.352		
+	0.0063	112.396		
+	0.0064	112.526		
+	0.0065	112.483		
+	0.0066	112.29		
+	0.0067	111.867		
+	0.0068	111.369		
+	0.0069	110.256		
+	0.007	108.626		
+	0.0071	106.511		
+	0.0072	103.246		
+	0.0073	98.587		
+	0.0074	91.962		
+	0.0075	82.29		
+	0.0076	73.42		
+	0.0077	66.384		
+	0.0078	60.145		
+	0.0079	54.112		
+	0.008	48.576		
+	0.0081	43.494		
+	0.0082	38.692		
+	0.0083	34.089		
+	0.0084	30.058		
+	0.0085	26.326		
+	0.0086	22.625		
+	0.0087	19.309		
+	0.0088	16.33		
+	0.0089	13.468		
+	0.009	10.738		
+	0.0091	8.498		
+	0.0092	6.365		
+	0.0093	4.399		
+	0.0094	2.782		
+	0.0095	1.407		
+	0.0096	0.194		
+	0.0097	-0.757		
+	0.0098	-1.46		
+	0.0099	-2.064		
+	0.01	-2.599		
+	0.0101	-2.804		
+	0.0102	-2.99		
+	0.0103	-3.158		
+	0.0104	-3.127		
+	0.0105	-2.99		
+	0.0106	-3.127		
+	0.0107	-3.077		
+	0.0108	-2.922		
+	0.0109	-2.941		
+	0.011	-2.947		
+	0.0111	-2.866		
+	0.0112	-2.791		
+	0.0113	-2.866		
+	0.0114	-2.717		
+	0.0115	-2.623		
+	0.0116	-2.655		
+	0.0117	-2.636		
+	0.0118	-2.431		
+	0.0119	-2.381		
+	0.012	-2.381		
+	0.0121	-2.269		
+	0.0122	-2.132		
+	0.0123	-2.138		
+	0.0124	-2.182		
+	0.0125	-2.057		
+	0.0126	-2.076		
+	0.0127	-2.207		
+	0.0128	-2.076		
+	0.0129	-2.032		
+	0.013	-2.032		
+	0.0131	-1.952		
+	0.0132	-1.952		
+	0.0133	-2.02		
+	0.0134	-1.914		
+	0.0135	-1.678		
+	0.0136	-1.703		
+	0.0137	-1.585		
+	0.0138	-1.529		
+	0.0139	-1.442		
+	0.014	-1.442		
+	0.0141	-1.336		
+	0.0142	-1.205		
+	0.0143	-1.274		
+	0.0144	-1.23		
+	0.0145	-1.081		
+	0.0146	-1.131		
+	0.0147	-1.081		
+	0.0148	-1.019		
+	0.0149	-0.931		
+	0.015	-0.963		
+	0.0151	-0.857		
+	0.0152	-0.72		
+	0.0153	-0.72		
+	0.0154	-0.676		
+	0.0155	-0.515		
+	0.0156	-0.521		
+	0.0157	-0.589		
+	0.0158	-0.471		
+	0.0159	-0.477		
+	0.016	-0.496		
+	0.0161	-0.372		
+	0.0162	-0.079		
+	0.0163	0.188		
+	0.0164	0.841		
+	0.0165	1.924		
+	0.0166	3.292		
+	0.0167	5.382		
+	0.0168	8.393		
+	0.0169	11.633		
+	0.017	15.366		
+	0.0171	19.515		
+	0.0172	24.118		
+	0.0173	28.926		
+	0.0174	34.114		
+	0.0175	39.743		
+	0.0176	45.77		
+	0.0177	51.879		
+	0.0178	58.385		
+	0.0179	64.979		
+	0.018	71.616		
+	0.0181	78.122		
+	0.0182	84.429		
+	0.0183	89.605		
+	0.0184	93.722		
+	0.0185	96.721		
+	0.0186	98.929		
+	0.0187	100.403		
+	0.0188	101.367		
+	0.0189	102.058		
+	0.019	102.58		
+	0.0191	103.04		
+	0.0192	103.575		
+	0.0193	104.073		
+	0.0194	104.739		
+	0.0195	105.553		
+	0.0196	106.3		
+	0.0197	107.084		
+	0.0198	107.843		
+	0.0199	108.589		
+	0.02	109.074		
+	0.0201	109.646		
+	0.0202	110.256		
+	0.0203	110.573		
+	0.0204	110.841		
+	0.0205	111.164		
+	0.0206	111.394		
+	0.0207	111.432		
+	0.0208	111.624		
+	0.0209	111.705		
+	0.021	111.712		
+	0.0211	111.705		
+	0.0212	111.805		
+	0.0213	111.755		
+	0.0214	111.755		
+	0.0215	111.792		
+	0.0216	111.712		
+	0.0217	111.587		
+	0.0218	111.593		
+	0.0219	111.792		
+	0.022	111.799		
+	0.0221	111.935		
+	0.0222	112.103		
+	0.0223	112.309		
+	0.0224	112.421		
+	0.0225	112.595		
+	0.0226	112.613		
+	0.0227	112.539		
+	0.0228	112.358		
+	0.0229	111.979		
+	0.023	111.276		
+	0.0231	110.206		
+	0.0232	108.626		
+	0.0233	106.325		
+	0.0234	103.04		
+	0.0235	98.531		
+	0.0236	91.937		
+	0.0237	82.171		
+	0.0238	73.488		
+	0.0239	66.54		
+	0.024	60.201		
+	0.0241	54.199		
+	0.0242	48.744		
+	0.0243	43.618		
+	0.0244	38.766		
+	0.0245	34.325		
+	0.0246	30.12		
+	0.0247	26.338		
+	0.0248	22.643		
+	0.0249	19.353		
+	0.025	16.205		
+	0.0251	13.363		
+	0.0252	10.844		
+	0.0253	8.573		
+	0.0254	6.415		
+	0.0255	4.598		
+	0.0256	3.012		
+	0.0257	1.55		
+	0.0258	0.381		
+	0.0259	-0.533		
+	0.026	-1.342		
+	0.0261	-2.032		
+	0.0262	-2.431		
+	0.0263	-2.779		
+	0.0264	-3.028		
+	0.0265	-3.14		
+	0.0266	-3.196		
+	0.0267	-3.165		
+	0.0268	-3.165		
+	0.0269	-3.046		
+	0.027	-2.941		
+	0.0271	-2.934		
+	0.0272	-2.922		
+	0.0273	-2.785		
+	0.0274	-2.729		
+	0.0275	-2.692		
+	0.0276	-2.58		
+	0.0277	-2.605		
+	0.0278	-2.536		
+	0.0279	-2.518		
+	0.028	-2.418		
+	0.0281	-2.443		
+	0.0282	-2.362		
+	0.0283	-2.35		
+	0.0284	-2.263		
+	0.0285	-2.25		
+	0.0286	-2.126		
+	0.0287	-2.126		
+	0.0288	-2.12		
+	0.0289	-2.064		
+	0.029	-1.995		
+	0.0291	-2.001		
+	0.0292	-1.933		
+	0.0293	-1.833		
+	0.0294	-1.921		
+	0.0295	-1.883		
+	0.0296	-1.765		
+	0.0297	-1.734		
+	0.0298	-1.753		
+	0.0299	-1.653		
+	0.03	-1.554		
+	0.0301	-1.628		
+	0.0302	-1.485		
+	0.0303	-1.323		
+	0.0304	-1.323		
+	0.0305	-1.298		
+	0.0306	-1.143		
+	0.0307	-0.994		
+	0.0308	-1.037		
+	0.0309	-0.9		
+	0.031	-0.876		
+	0.0311	-0.9		
+	0.0312	-0.9		
+	0.0313	-0.77		
+	0.0314	-0.788		
+	0.0315	-0.77		
+	0.0316	-0.714		
+	0.0317	-0.62		
+	0.0318	-0.701		
+	0.0319	-0.546		
+	0.032	-0.49		
+	0.0321	-0.459		
+	0.0322	-0.428		
+	0.0323	-0.272		
+	0.0324	-0.067		
+	0.0325	0.313		
+	0.0326	0.966		
+	0.0327	1.893		
+	0.0328	3.217		
+	0.0329	5.233		
+	0.033	8.163		
+	0.0331	11.31		
+	0.0332	14.974		
+	0.0333	19.085		
+	0.0334	23.496		
+	0.0335	28.248		
+	0.0336	33.535		
+	0.0337	39.04		
+	0.0338	44.937		
+	0.0339	51.12		
+	0.034	57.651		
+	0.0341	64.182		
+	0.0342	70.745		
+	0.0343	77.289		
+	0.0344	83.552		
+	0.0345	88.821		
+	0.0346	93.057		
+	0.0347	96.223		
+	0.0348	98.413		
+	0.0349	99.961		
+	0.035	101.069		
+	0.0351	101.703		
+	0.0352	102.25		
+	0.0353	102.823		
+	0.0354	103.37		
+	0.0355	103.886		
+	0.0356	104.602		
+	0.0357	105.466		
+	0.0358	106.144		
+	0.0359	106.941		
+	0.036	107.737		
+	0.0361	108.353		
+	0.0362	108.937		
+	0.0363	109.578		
+	0.0364	110.094		
+	0.0365	110.331		
+	0.0366	110.648		
+	0.0367	110.953		
+	0.0368	111.096		
+	0.0369	111.351		
+	0.037	111.5		
+	0.0371	111.649		
+	0.0372	111.662		
+	0.0373	111.712		
+	0.0374	111.768		
+	0.0375	111.755		
+	0.0376	111.805		
+	0.0377	111.768		
+	0.0378	111.687		
+	0.0379	111.55		
+	0.038	111.693		
+	0.0381	111.593		
+	0.0382	111.612		
+	0.0383	111.768		
+	0.0384	111.985		
+	0.0385	112.097		
+	0.0386	112.296		
+	0.0387	112.489		
+	0.0388	112.526		
+	0.0389	112.502		
+	0.039	112.402		
+	0.0391	112.147		
+	0.0392	111.376		
+	0.0393	110.455		
+	0.0394	108.987		
+	0.0395	106.623		
+	0.0396	103.607		
+	0.0397	99.377		
+	0.0398	93.113		
+	0.0399	83.615		
+	0.04	74.744		
+	0.0401	67.572		
+	0.0402	61.141		
+	0.0403	55.194		
+	0.0404	49.789		
+	0.0405	44.489		
+	0.0406	39.631		
+	0.0407	35.277		
+	0.0408	31.003		
+	0.0409	27.035		
+	0.041	23.502		
+	0.0411	20.012		
+	0.0412	16.809		
+	0.0413	13.935		
+	0.0414	11.341		
+	0.0415	8.828		
+	0.0416	6.701		
+	0.0417	4.884		
+	0.0418	3.168		
+	0.0419	1.749		
+	0.042	0.611		
+	0.0421	-0.328		
+	0.0422	-1.311		
+	0.0423	-1.765		
+	0.0424	-2.219		
+	0.0425	-2.642		
+	0.0426	-2.872		
+	0.0427	-2.934		
+	0.0428	-3.152		
+	0.0429	-3.239		
+	0.043	-3.096		
+	0.0431	-3.04		
+	0.0432	-3.146		
+	0.0433	-2.997		
+	0.0434	-2.953		
+	0.0435	-2.947		
+	0.0436	-2.866		
+	0.0437	-2.655		
+	0.0438	-2.592		
+	0.0439	-2.648		
+	0.044	-2.368		
+	0.0441	-2.362		
+	0.0442	-2.393		
+	0.0443	-2.343		
+	0.0444	-2.232		
+	0.0445	-2.331		
+	0.0446	-2.3		
+	0.0447	-2.163		
+	0.0448	-2.188		
+	0.0449	-2.294		
+	0.045	-2.2		
+	0.0451	-2.082		
+	0.0452	-2.107		
+	0.0453	-2.001		
+	0.0454	-1.852		
+	0.0455	-1.939		
+	0.0456	-1.883		
+	0.0457	-1.715		
+	0.0458	-1.672		
+	0.0459	-1.784		
+	0.046	-1.585		
+	0.0461	-1.566		
+	0.0462	-1.585		
+	0.0463	-1.572		
+	0.0464	-1.354		
+	0.0465	-1.448		
+	0.0466	-1.473		
+	0.0467	-1.23		
+	0.0468	-1.131		
+	0.0469	-1.187		
+	0.047	-0.963		
+	0.0471	-0.801		
+	0.0472	-0.931		
+	0.0473	-0.838		
+	0.0474	-0.664		
+	0.0475	-0.708		
+	0.0476	-0.745		
+	0.0477	-0.627		
+	0.0478	-0.62		
+	0.0479	-0.708		
+	0.048	-0.571		
+	0.0481	-0.552		
+	0.0482	-0.645		
+	0.0483	-0.67		
+	0.0484	-0.465		
+	0.0485	-0.39		
+	0.0486	-0.21		
+	0.0487	0.356		
+	0.0488	0.991		
+	0.0489	1.861		
+	0.049	3.242		
+	0.0491	5.301		
+	0.0492	8.026		
+	0.0493	11.173		
+	0.0494	14.787		
+	0.0495	18.743		
+	0.0496	23.066		
+	0.0497	27.887		
+	0.0498	33		
+	0.0499	38.343		
+	0.05	44.203		
+	0.0501	50.454		
+	0.0502	56.718		
+	0.0503	63.224		
+	0.0504	69.924		
+	0.0505	76.306		
+	0.0506	82.563		
+	0.0507	88.174		
+	0.0508	92.522		
+	0.0509	95.682		
+	0.051	98.046		
+	0.0511	99.793		
+	0.0512	100.764		
+	0.0513	101.386		
+	0.0514	102.126		
+	0.0515	102.543		
+	0.0516	102.96		
+	0.0517	103.656		
+	0.0518	104.353		
+	0.0519	104.963		
+	0.052	105.889		
+	0.0521	106.841		
+	0.0522	107.476		
+	0.0523	108.185		
+	0.0524	108.869		
+	0.0525	109.435		
+	0.0526	109.827		
+	0.0527	110.268		
+	0.0528	110.648		
+	0.0529	110.754		
+	0.053	111.04		
+	0.0531	111.295		
+	0.0532	111.301		
+	0.0533	111.295		
+	0.0534	111.562		
+	0.0535	111.568		
+	0.0536	111.519		
+	0.0537	111.755		
+	0.0538	111.73		
+	0.0539	111.643		
+	0.054	111.624		
+	0.0541	111.656		
+	0.0542	111.531		
+	0.0543	111.581		
+	0.0544	111.631		
+	0.0545	111.743		
+	0.0546	111.736		
+	0.0547	112.035		
+	0.0548	112.159		
+	0.0549	112.246		
+	0.055	112.246		
+	0.0551	112.377		
+	0.0552	112.222		
+	0.0553	111.898		
+	0.0554	111.425		
+	0.0555	110.536		
+	0.0556	108.968		
+	0.0557	107.028		
+	0.0558	104.135		
+	0.0559	99.974		
+	0.056	94.121		
+	0.0561	85.182		
+	0.0562	75.814		
+	0.0563	68.418		
+	0.0564	62.123		
+	0.0565	56.046		
+	0.0566	50.38		
+	0.0567	45.223		
+	0.0568	40.371		
+	0.0569	35.737		
+	0.057	31.601		
+	0.0571	27.806		
+	0.0572	23.981		
+	0.0573	20.497		
+	0.0574	17.499		
+	0.0575	14.569		
+	0.0576	11.783		
+	0.0577	9.357		
+	0.0578	7.242		
+	0.0579	5.146		
+	0.058	3.441		
+	0.0581	2.06		
+	0.0582	0.754		
+	0.0583	-0.39		
+	0.0584	-1.131		
+	0.0585	-1.765		
+	0.0586	-2.3		
+	0.0587	-2.561		
+	0.0588	-2.692		
+	0.0589	-2.978		
+	0.059	-3.09		
+	0.0591	-2.941		
+	0.0592	-2.978		
+	0.0593	-3.084		
+	0.0594	-2.953		
+	0.0595	-2.966		
+	0.0596	-3.077		
+	0.0597	-2.941		
+	0.0598	-2.822		
+	0.0599	-2.835		
+	0.06	-2.754		
+	0.0601	-2.561		
+	0.0602	-2.474		
+	0.0603	-2.53		
+	0.0604	-2.35		
+	0.0605	-2.269		
+	0.0606	-2.325		
+	0.0607	-2.232		
+	0.0608	-2.057		
+	0.0609	-2.163		
+	0.061	-2.225		
+	0.0611	-2.088		
+	0.0612	-2.157		
+	0.0613	-2.194		
+	0.0614	-2.07		
+	0.0615	-2.001		
+	0.0616	-2.07		
+	0.0617	-2.001		
+	0.0618	-1.871		
+	0.0619	-1.846		
+	0.062	-1.784		
+	0.0621	-1.622		
+	0.0622	-1.597		
+	0.0623	-1.622		
+	0.0624	-1.442		
+	0.0625	-1.33		
+	0.0626	-1.423		
+	0.0627	-1.361		
+	0.0628	-1.211		
+	0.0629	-1.298		
+	0.063	-1.236		
+	0.0631	-1.062		
+	0.0632	-1.106		
+	0.0633	-1.099		
+	0.0634	-0.907		
+	0.0635	-0.869		
+	0.0636	-0.813		
+	0.0637	-0.745		
+	0.0638	-0.589		
+	0.0639	-0.645		
+	0.064	-0.583		
+	0.0641	-0.484		
+	0.0642	-0.515		
+	0.0643	-0.564		
+	0.0644	-0.54		
+	0.0645	-0.515		
+	0.0646	-0.577		
+	0.0647	-0.446		
+	0.0648	-0.21		
+	0.0649	0.138		
+	0.065	0.68		
+	0.0651	1.756		
+	0.0652	3.043		
+	0.0653	5.015		
+	0.0654	7.764		
+	0.0655	10.993		
+	0.0656	14.489		
+	0.0657	18.382		
+	0.0658	22.855		
+	0.0659	27.47		
+	0.066	32.409		
+	0.0661	37.864		
+	0.0662	43.593		
+	0.0663	49.565		
+	0.0664	55.866		
+	0.0665	62.347		
+	0.0666	68.767		
+	0.0667	75.192		
+	0.0668	81.593		
+	0.0669	87.241		
+	0.067	91.657		
+	0.0671	95.097		
+	0.0672	97.647		
+	0.0673	99.283		
+	0.0674	100.527		
+	0.0675	101.436		
+	0.0676	101.89		
+	0.0677	102.195		
+	0.0678	102.854		
+	0.0679	103.289		
+	0.068	103.974		
+	0.0681	104.72		
+	0.0682	105.516		
+	0.0683	106.219		
+	0.0684	107.009		
+	0.0685	107.874		
+	0.0686	108.508		
+	0.0687	109.037		
+	0.0688	109.721		
+	0.0689	110.001		
+	0.069	110.3		
+	0.0691	110.679		
+	0.0692	110.934		
+	0.0693	111.027		
+	0.0694	111.108		
+	0.0695	111.22		
+	0.0696	111.195		
+	0.0697	111.214		
+	0.0698	111.481		
+	0.0699	111.444		
+	0.07	111.351		
+	0.0701	111.438		
+	0.0702	111.537		
+	0.0703	111.413		
+	0.0704	111.444		
+	0.0705	111.525		
+	0.0706	111.575		
+	0.0707	111.581		
+	0.0708	111.824		
+	0.0709	111.991		
+	0.071	111.923		
+	0.0711	112.147		
+	0.0712	112.24		
+	0.0713	112.159		
+	0.0714	112.01		
+	0.0715	111.805		
+	0.0716	111.295		
+	0.0717	110.287		
+	0.0718	109.093		
+	0.0719	107.202		
+	0.072	104.378		
+	0.0721	100.627		
+	0.0722	95.209		
+	0.0723	86.712		
+	0.0724	77.201		
+	0.0725	69.768		
+	0.0726	63.113		
+	0.0727	56.948		
+	0.0728	51.35		
+	0.0729	46.088		
+	0.073	41.093		
+	0.0731	36.508		
+	0.0732	32.26		
+	0.0733	28.173		
+	0.0734	24.553		
+	0.0735	21.132		
+	0.0736	17.891		
+	0.0737	14.856		
+	0.0738	12.318		
+	0.0739	9.786		
+	0.074	7.441		
+	0.0741	5.513		
+	0.0742	3.759		
+	0.0743	2.16		
+	0.0744	0.866		
+	0.0745	-0.117		
+	0.0746	-1.093		
+	0.0747	-1.852		
+	0.0748	-2.269		
+	0.0749	-2.661		
+	0.075	-2.978		
+	0.0751	-3.152		
+	0.0752	-3.046		
+	0.0753	-3.146		
+	0.0754	-3.165		
+	0.0755	-3.071		
+	0.0756	-2.984		
+	0.0757	-2.966		
+	0.0758	-2.934		
+	0.0759	-2.829		
+	0.076	-2.885		
+	0.0761	-2.804		
+	0.0762	-2.723		
+	0.0763	-2.748		
+	0.0764	-2.686		
+	0.0765	-2.655		
+	0.0766	-2.511		
+	0.0767	-2.543		
+	0.0768	-2.443		
+	0.0769	-2.306		
+	0.077	-2.288		
+	0.0771	-2.238		
+	0.0772	-2.144		
+	0.0773	-2.07		
+	0.0774	-2.12		
+	0.0775	-2.039		
+	0.0776	-1.995		
+	0.0777	-2.051		
+	0.0778	-2.113		
+	0.0779	-1.983		
+	0.078	-1.97		
+	0.0781	-1.952		
+	0.0782	-1.865		
+	0.0783	-1.865		
+	0.0784	-1.84		
+	0.0785	-1.678		
+	0.0786	-1.56		
+	0.0787	-1.56		
+	0.0788	-1.379		
+	0.0789	-1.255		
+	0.079	-1.305		
+	0.0791	-1.205		
+	0.0792	-1.087		
+	0.0793	-1.081		
+	0.0794	-1.112		
+	0.0795	-1.075		
+	0.0796	-1		
+	0.0797	-0.907		
+	0.0798	-0.907		
+	0.0799	-0.813		
+	0.08	-0.77		
+	0.0801	-0.751		
+	0.0802	-0.633		
+	0.0803	-0.564		
+	0.0804	-0.515		
+	0.0805	-0.515		
+	0.0806	-0.465		
+	0.0807	-0.533		
+	0.0808	-0.428		
+	0.0809	-0.316		
+	0.081	-0.086		
+	0.0811	0.132		
+	0.0812	0.742		
+	0.0813	1.494		
+	0.0814	2.72		
+	0.0815	4.536		
+	0.0816	7.23		
+	0.0817	10.253		
+	0.0818	13.736		
+	0.0819	17.667		
+	0.082	21.99		
+	0.0821	26.593		
+	0.0822	31.545		
+	0.0823	36.819		
+	0.0824	42.399		
+	0.0825	48.476		
+	0.0826	54.721		
+	0.0827	61.072		
+	0.0828	67.373		
+	0.0829	73.867		
+	0.083	80.156		
+	0.0831	85.879		
+	0.0832	90.563		
+	0.0833	94.195		
+	0.0834	96.783		
+	0.0835	98.78		
+	0.0836	100.148		
+	0.0837	101.075		
+	0.0838	101.703		
+	0.0839	102.201		
+	0.084	102.748		
+	0.0841	103.215		
+	0.0842	103.83		
+	0.0843	104.633		
+	0.0844	105.274		
+	0.0845	106.057		
+	0.0846	106.847		
+	0.0847	107.612		
+	0.0848	108.166		
+	0.0849	108.869		
+	0.085	109.373		
+	0.0851	109.777		
+	0.0852	110.181		
+	0.0853	110.542		
+	0.0854	110.828		
+	0.0855	110.928		
+	0.0856	111.164		
+	0.0857	111.307		
+	0.0858	111.301		
+	0.0859	111.413		
+	0.086	111.444		
+	0.0861	111.382		
+	0.0862	111.407		
+	0.0863	111.457		
+	0.0864	111.413		
+	0.0865	111.32		
+	0.0866	111.369		
+	0.0867	111.32		
+	0.0868	111.394		
+	0.0869	111.612		
+	0.087	111.743		
+	0.0871	111.886		
+	0.0872	112.023		
+	0.0873	112.215		
+	0.0874	112.315		
+	0.0875	112.321		
+	0.0876	112.315		
+	0.0877	112.023		
+	0.0878	111.5		
+	0.0879	110.741		
+	0.088	109.566		
+	0.0881	107.755		
+	0.0882	105.249		
+	0.0883	101.896		
+	0.0884	96.951		
+	0.0885	89.735		
+	0.0886	80.088		
+	0.0887	72.02		
+	0.0888	65.271		
+	0.0889	59.069		
+	0.089	53.347		
+	0.0891	47.941		
+	0.0892	42.946		
+	0.0893	38.25		
+	0.0894	33.815		
+	0.0895	29.679		
+	0.0896	25.859		
+	0.0897	22.314		
+	0.0898	18.992		
+	0.0899	15.95		
+	0.09	13.164		
+	0.0901	10.632		
+	0.0902	8.256		
+	0.0903	6.247		
+	0.0904	4.48		
+	0.0905	2.732		
+	0.0906	1.426		
+	0.0907	0.4		
+	0.0908	-0.676		
+	0.0909	-1.386		
+	0.091	-1.933		
+	0.0911	-2.493		
+	0.0912	-2.785		
+	0.0913	-3.015		
+	0.0914	-3.084		
+	0.0915	-3.27		
+	0.0916	-3.221		
+	0.0917	-3.152		
+	0.0918	-3.127		
+	0.0919	-3.028		
+	0.092	-2.866		
+	0.0921	-2.841		
+	0.0922	-2.872		
+	0.0923	-2.729		
+	0.0924	-2.648		
+	0.0925	-2.623		
+	0.0926	-2.505		
+	0.0927	-2.48		
+	0.0928	-2.499		
+	0.0929	-2.524		
+	0.093	-2.387		
+	0.0931	-2.375		
+	0.0932	-2.368		
+	0.0933	-2.275		
+	0.0934	-2.163		
+	0.0935	-2.219		
+	0.0936	-2.101		
+	0.0937	-2.008		
+	0.0938	-2.032		
+	0.0939	-2.076		
+	0.094	-1.914		
+	0.0941	-1.896		
+	0.0942	-1.939		
+	0.0943	-1.746		
+	0.0944	-1.809		
+	0.0945	-1.865		
+	0.0946	-1.802		
+	0.0947	-1.634		
+	0.0948	-1.684		
+	0.0949	-1.616		
+	0.095	-1.454		
+	0.0951	-1.41		
+	0.0952	-1.404		
+	0.0953	-1.224		
+	0.0954	-1.143		
+	0.0955	-1.168		
+	0.0956	-1.037		
+	0.0957	-0.863		
+	0.0958	-0.826		
+	0.0959	-0.876		
+	0.096	-0.739		
+	0.0961	-0.708		
+	0.0962	-0.832		
+	0.0963	-0.757		
+	0.0964	-0.639		
+	0.0965	-0.757		
+	0.0966	-0.664		
+	0.0967	-0.577		
+	0.0968	-0.596		
+	0.0969	-0.558		
+	0.097	-0.39		
+	0.0971	-0.322		
+	0.0972	-0.278		
+	0.0973	0.132		
+	0.0974	0.667		
+	0.0975	1.239		
+	0.0976	2.303		
+	0.0977	3.895		
+	0.0978	6.178		
+	0.0979	9.002		
+	0.098	12.311		
+	0.0981	16.044		
+	0.0982	20.074		
+	0.0983	24.541		
+	0.0984	29.374		
+	0.0985	34.449		
+	0.0986	40.029		
+	0.0987	45.926		
+	0.0988	52.034		
+	0.0989	58.298		
+	0.099	64.711		
+	0.0991	71.149		
+	0.0992	77.425		
+	0.0993	83.434		
+	0.0994	88.647		
+	0.0995	92.584		
+	0.0996	95.595		
+	0.0997	97.94		
+	0.0998	99.538		
+	0.0999	100.459		
+	0.1	101.274		
+	0.1001	101.884		
+	0.1002	102.269		
+	0.1003	102.947		
+	0.1004	103.588		
+	0.1005	104.166		
+	0.1006	104.969		
+	0.1007	105.883		
+	0.1008	106.574		
+	0.1009	107.258		
+	0.101	107.998		
+	0.1011	108.707		
+	0.1012	109.13		
+	0.1013	109.547		
+	0.1014	110.113		
+	0.1015	110.312		
+	0.1016	110.53		
+	0.1017	110.872		
+	0.1018	111.052		
+	0.1019	111.108		
+	0.102	111.282		
+	0.1021	111.438		
+	0.1022	111.401		
+	0.1023	111.494		
+	0.1024	111.637		
+	0.1025	111.593		
+	0.1026	111.575		
+	0.1027	111.6		
+	0.1028	111.575		
+	0.1029	111.444		
+	0.103	111.587		
+	0.1031	111.68		
+	0.1032	111.699		
+	0.1033	111.824		
+	0.1034	112.159		
+	0.1035	112.166		
+	0.1036	112.302		
+	0.1037	112.489		
+	0.1038	112.47		
+	0.1039	112.278		
+	0.104	112.085		
+	0.1041	111.606		
+	0.1042	110.505		
+	0.1043	109.012		
+	0.1044	107.077		
+	0.1045	104.061		
+	0.1046	99.986		
+	0.1047	94.481		
+	0.1048	85.636		
+	0.1049	76.374		
+	0.105	69.059		
+	0.1051	62.752		
+	0.1052	56.612		
+	0.1053	51.101		
+	0.1054	45.988		
+	0.1055	41.099		
+	0.1056	36.428		
+	0.1057	32.303		
+	0.1058	28.36		
+	0.1059	24.553		
+	0.106	21.151		
+	0.1061	18.034		
+	0.1062	14.893		
+	0.1063	12.125		
+	0.1064	9.798		
+	0.1065	7.466		
+	0.1066	5.457		
+	0.1067	3.808		
+	0.1068	2.235		
+	0.1069	0.866		
+	0.107	-0.073		
+	0.1071	-0.838		
+	0.1072	-1.622		
+	0.1073	-2.176		
+	0.1074	-2.431		
+	0.1075	-2.729		
+	0.1076	-3.009		
+	0.1077	-2.99		
+	0.1078	-3.059		
+	0.1079	-3.165		
+	0.108	-3.14		
+	0.1081	-2.966		
+	0.1082	-3.034		
+	0.1083	-3.003		
+	0.1084	-2.903		
+	0.1085	-2.866		
+	0.1086	-2.76		
+	0.1087	-2.679		
+	0.1088	-2.493		
+	0.1089	-2.561		
+	0.109	-2.474		
+	0.1091	-2.275		
+	0.1092	-2.356		
+	0.1093	-2.387		
+	0.1094	-2.232		
+	0.1095	-2.225		
+	0.1096	-2.325		
+	0.1097	-2.132		
+	0.1098	-2.132		
+	0.1099	-2.207		
+	0.11	-2.151		
+	0.1101	-2.039		
+	0.1102	-2.051		
+	0.1103	-2.045		
+	0.1104	-1.815		
+	0.1105	-1.815		
+	0.1106	-1.858		
+	0.1107	-1.697		
+	0.1108	-1.634		
+	0.1109	-1.665		
+	0.111	-1.554		
+	0.1111	-1.485		
+	0.1112	-1.473		
+	0.1113	-1.554		
+	0.1114	-1.354		
+	0.1115	-1.292		
+	0.1116	-1.317		
+	0.1117	-1.118		
+	0.1118	-1.087		
+	0.1119	-1.019		
+	0.112	-0.95		
+	0.1121	-0.776		
+	0.1122	-0.82		
+	0.1123	-0.826		
+	0.1124	-0.639		
+	0.1125	-0.552		
+	0.1126	-0.701		
+	0.1127	-0.62		
+	0.1128	-0.502		
+	0.1129	-0.664		
+	0.113	-0.602		
+	0.1131	-0.428		
+	0.1132	-0.49		
+	0.1133	-0.54		
+	0.1134	-0.328		
+	0.1135	-0.129		
+	0.1136	0.219		
+	0.1137	0.922		
+	0.1138	1.868		
+	0.1139	3.012		
+	0.114	4.972		
+	0.1141	7.814		
+	0.1142	10.949		
+	0.1143	14.314		
+	0.1144	18.271		
+	0.1145	22.494		
+	0.1146	26.985		
+	0.1147	32.073		
+	0.1148	37.392		
+	0.1149	42.897		
+	0.115	48.881		
+	0.1151	55.169		
+	0.1152	61.433		
+	0.1153	67.747		
+	0.1154	74.259		
+	0.1155	80.492		
+	0.1156	86.034		
+	0.1157	90.712		
+	0.1158	94.388		
+	0.1159	96.895		
+	0.116	98.761		
+	0.1161	100.167		
+	0.1162	101.013		
+	0.1163	101.597		
+	0.1164	102.157		
+	0.1165	102.686		
+	0.1166	103.096		
+	0.1167	103.762		
+	0.1168	104.62		
+	0.1169	105.342		
+	0.117	106.151		
+	0.1171	107.109		
+	0.1172	107.724		
+	0.1173	108.433		
+	0.1174	109.062		
+	0.1175	109.634		
+	0.1176	109.945		
+	0.1177	110.318		
+	0.1178	110.685		
+	0.1179	110.822		
+	0.118	110.99		
+	0.1181	111.307		
+	0.1182	111.382		
+	0.1183	111.338		
+	0.1184	111.556		
+	0.1185	111.693		
+	0.1186	111.643		
+	0.1187	111.755		
+	0.1188	111.898		
+	0.1189	111.792		
+	0.119	111.824		
+	0.1191	111.935		
+	0.1192	111.96		
+	0.1193	111.911		
+	0.1194	112.029		
+	0.1195	112.147		
+	0.1196	112.178		
+	0.1197	112.377		
+	0.1198	112.62		
+	0.1199	112.626		
+	0.12	112.607		
+	0.1201	112.701		
+	0.1202	112.557		
+	0.1203	111.998		
+	0.1204	111.519		
+	0.1205	110.48		
+	0.1206	108.676		
+	0.1207	106.412		
+	0.1208	103.314		
+	0.1209	98.68		
+	0.121	92.062		
+	0.1211	82.551		
+	0.1212	74.01		
+	0.1213	67.031		
+	0.1214	60.823		
+	0.1215	55.07		
+	0.1216	49.459		
+	0.1217	44.346		
+	0.1218	39.737		
+	0.1219	35.277		
+	0.122	31.115		
+	0.1221	27.383		
+	0.1222	23.726		
+	0.1223	20.249		
+	0.1224	17.188		
+	0.1225	14.445		
+	0.1226	11.665		
+	0.1227	9.12		
+	0.1228	7.136		
+	0.1229	5.115		
+	0.123	3.354		
+	0.1231	1.924		
+	0.1232	0.742		
+	0.1233	-0.421		
+	0.1234	-1.205		
+	0.1235	-1.734		
+	0.1236	-2.238		
+	0.1237	-2.661		
+	0.1238	-2.686		
+	0.1239	-2.903		
+	0.124	-3.084		
+	0.1241	-3.015		
+	0.1242	-2.885		
+	0.1243	-3.015		
+	0.1244	-2.99		
+	0.1245	-2.928		
+	0.1246	-2.953		
+	0.1247	-2.816		
+	0.1248	-2.742		
+	0.1249	-2.791		
+	0.125	-2.698		
+	0.1251	-2.599		
+	0.1252	-2.418		
+	0.1253	-2.468		
+	0.1254	-2.368		
+	0.1255	-2.194		
+	0.1256	-2.244		
+	0.1257	-2.238		
+	0.1258	-2.076		
+	0.1259	-2.126		
+	0.126	-2.107		
+	0.1261	-2.07		
+	0.1262	-1.989		
+	0.1263	-2.151		
+	0.1264	-2.014		
+	0.1265	-1.958		
+	0.1266	-2.001		
+	0.1267	-2.001		
+	0.1268	-1.833		
+	0.1269	-1.74		
+	0.127	-1.74		
+	0.1271	-1.572		
+	0.1272	-1.541		
+	0.1273	-1.554		
+	0.1274	-1.435		
+	0.1275	-1.342		
+	0.1276	-1.267		
+	0.1277	-1.286		
+	0.1278	-1.199		
+	0.1279	-1.099		
+	0.128	-1.193		
+	0.1281	-1.056		
+	0.1282	-0.969		
+	0.1283	-0.981		
+	0.1284	-0.876		
+	0.1285	-0.726		
+	0.1286	-0.701		
+	0.1287	-0.683		
+	0.1288	-0.564		
+	0.1289	-0.515		
+	0.129	-0.54		
+	0.1291	-0.533		
+	0.1292	-0.421		
+	0.1293	-0.434		
+	0.1294	-0.527		
+	0.1295	-0.378		
+	0.1296	-0.334		
+	0.1297	-0.316		
+	0.1298	0.02		
+	0.1299	0.393		
+	0.13	0.991		
+	0.1301	1.936		
+	0.1302	3.553		
+	0.1303	5.587		
+	0.1304	8.424		
+	0.1305	11.665		
+	0.1306	15.21		
+	0.1307	19.154		
+	0.1308	23.545		
+	0.1309	28.229		
+	0.131	33.199		
+	0.1311	38.518		
+	0.1312	44.259		
+	0.1313	50.106		
+	0.1314	56.283		
+	0.1315	62.727		
+	0.1316	68.966		
+	0.1317	75.242		
+	0.1318	81.462		
+	0.1319	87.011		
+	0.132	91.508		
+	0.1321	94.942		
+	0.1322	97.43		
+	0.1323	99.296		
+	0.1324	100.478		
+	0.1325	101.473		
+	0.1326	102.07		
+	0.1327	102.437		
+	0.1328	103.016		
+	0.1329	103.582		
+	0.133	104.092		
+	0.1331	104.844		
+	0.1332	105.697		
+	0.1333	106.468		
+	0.1334	107.245		
+	0.1335	108.017		
+	0.1336	108.794		
+	0.1337	109.304		
+	0.1338	109.883		
+	0.1339	110.356		
+	0.134	110.648		
+	0.1341	110.953		
+	0.1342	111.332		
+	0.1343	111.519		
+	0.1344	111.531		
+	0.1345	111.774		
+	0.1346	111.848		
+	0.1347	111.867		
+	0.1348	111.929		
+	0.1349	112.035		
+	0.135	111.96		
+	0.1351	112.023		
+	0.1352	112.116		
+	0.1353	112.141		
+	0.1354	112.191		
+	0.1355	112.271		
+	0.1356	112.327		
+	0.1357	112.433		
+	0.1358	112.613		
+	0.1359	112.781		
+	0.136	112.875		
+	0.1361	112.999		
+	0.1362	113.161		
+	0.1363	113.18		
+	0.1364	113.08		
+	0.1365	113.012		
+	0.1366	112.533		
+	0.1367	111.861		
+	0.1368	110.803		
+	0.1369	109.143		
+	0.137	106.798		
+	0.1371	103.644		
+	0.1372	99.091		
+	0.1373	92.572		
+	0.1374	83.024		
+	0.1375	74.608		
+	0.1376	67.778		
+	0.1377	61.371		
+	0.1378	55.505		
+	0.1379	50.1		
+	0.138	44.999		
+	0.1381	40.234		
+	0.1382	35.756		
+	0.1383	31.613		
+	0.1384	27.688		
+	0.1385	24.049		
+	0.1386	20.728		
+	0.1387	17.543		
+	0.1388	14.663		
+	0.1389	12.056		
+	0.139	9.618		
+	0.1391	7.354		
+	0.1392	5.475		
+	0.1393	3.696		
+	0.1394	2.185		
+	0.1395	0.991		
+	0.1396	-0.104		
+	0.1397	-1.012		
+	0.1398	-1.709		
+	0.1399	-2.157		
+	0.14	-2.555		
+	0.1401	-2.86		
+	0.1402	-2.941		
+	0.1403	-2.934		
+	0.1404	-3.009		
+	0.1405	-2.978		
+	0.1406	-2.878		
+	0.1407	-2.829		
+	0.1408	-2.866		
+	0.1409	-2.742		
+	0.141	-2.735		
+	0.1411	-2.71		
+	0.1412	-2.642		
+	0.1413	-2.574		
+	0.1414	-2.555		
+	0.1415	-2.474		
+	0.1416	-2.487		
+	0.1417	-2.387		
+	0.1418	-2.393		
+	0.1419	-2.263		
+	0.142	-2.132		
+	0.1421	-2.151		
+	0.1422	-2.107		
+	0.1423	-2.02		
+	0.1424	-2.001		
+	0.1425	-1.958		
+	0.1426	-1.939		
+	0.1427	-1.933		
+	0.1428	-1.989		
+	0.1429	-1.939		
+	0.143	-1.858		
+	0.1431	-1.846		
+	0.1432	-1.74		
+	0.1433	-1.709		
+	0.1434	-1.647		
+	0.1435	-1.597		
+	0.1436	-1.498		
+	0.1437	-1.386		
+	0.1438	-1.342		
+	0.1439	-1.274		
+	0.144	-1.218		
+	0.1441	-1.174		
+	0.1442	-1.087		
+	0.1443	-0.975		
+	0.1444	-0.981		
+	0.1445	-0.931		
+	0.1446	-0.894		
+	0.1447	-0.788		
+	0.1448	-0.732		
+	0.1449	-0.695		
+	0.145	-0.676		
+	0.1451	-0.633		
+	0.1452	-0.533		
+	0.1453	-0.365		
+	0.1454	-0.434		
+	0.1455	-0.434		
+	0.1456	-0.328		
+	0.1457	-0.309		
+	0.1458	-0.272		
+	0.1459	-0.185		
+	0.146	-0.067		
+	0.1461	0.182		
+	0.1462	0.617		
+	0.1463	1.407		
+	0.1464	2.552		
+	0.1465	4.244		
+	0.1466	6.614		
+	0.1467	9.587		
+	0.1468	12.809		
+	0.1469	16.61		
+	0.147	20.765		
+	0.1471	25.194		
+	0.1472	29.94		
+	0.1473	35.103		
+	0.1474	40.508		
+	0.1475	46.243		
+	0.1476	52.333		
+	0.1477	58.59		
+	0.1478	64.736		
+	0.1479	71.006		
+	0.148	77.351		
+	0.1481	83.285		
+	0.1482	88.466		
+	0.1483	92.702		
+	0.1484	95.844		
+	0.1485	98.064		
+	0.1486	99.831		
+	0.1487	101		
+	0.1488	101.734		
+	0.1489	102.362		
+	0.149	102.916		
+	0.1491	103.345		
+	0.1492	103.936		
+	0.1493	104.614		
+	0.1494	105.373		
+	0.1495	106.039		
+	0.1496	106.816		
+	0.1497	107.78		
+	0.1498	108.384		
+	0.1499	109.062		
+	0.15	109.671		
+	0.1501	110.094		
+	0.1502	110.567		
+	0.1503	110.984		
+	0.1504	111.239		
+	0.1505	111.519		
+	0.1506	111.749		
+	0.1507	111.948		
+	0.1508	111.979		
+	0.1509	112.11		
+	0.151	112.191		
+	0.1511	112.191		
+	0.1512	112.271		
+	0.1513	112.296		
+	0.1514	112.365		
+	0.1515	112.346		
+	0.1516	112.278		
+	0.1517	112.421		
+	0.1518	112.396		
+	0.1519	112.489		
+	0.152	112.763		
+	0.1521	112.987		
+	0.1522	113.049		
+	0.1523	113.323		
+	0.1524	113.522		
+	0.1525	113.559		
+	0.1526	113.584		
+	0.1527	113.54		
+	0.1528	113.217		
+	0.1529	112.719		
+	0.153	111.985		
+	0.1531	110.754		
+	0.1532	108.944		
+	0.1533	106.487		
+	0.1534	103.04		
+	0.1535	98.195		
+	0.1536	91.035		
+	0.1537	81.556		
+	0.1538	73.444		
+	0.1539	66.745		
+	0.154	60.631		
+	0.1541	54.852		
+	0.1542	49.44		
+	0.1543	44.458		
+	0.1544	39.78		
+	0.1545	35.351		
+	0.1546	31.178		
+	0.1547	27.47		
+	0.1548	23.775		
+	0.1549	20.398		
+	0.155	17.269		
+	0.1551	14.402		
+	0.1552	11.652		
+	0.1553	9.382		
+	0.1554	7.267		
+	0.1555	5.27		
+	0.1556	3.547		
+	0.1557	2.172		
+	0.1558	0.891		
+	0.1559	-0.16		
+	0.156	-0.913		
+	0.1561	-1.572		
+	0.1562	-2.182		
+	0.1563	-2.499		
+	0.1564	-2.723		
+	0.1565	-2.922		
+	0.1566	-3.04		
+	0.1567	-2.997		
+	0.1568	-3.028		
+	0.1569	-3.015		
+	0.157	-2.86		
+	0.1571	-2.748		
+	0.1572	-2.735		
+	0.1573	-2.717		
+	0.1574	-2.574		
+	0.1575	-2.53		
+	0.1576	-2.561		
+	0.1577	-2.387		
+	0.1578	-2.362		
+	0.1579	-2.443		
+	0.158	-2.325		
+	0.1581	-2.232		
+	0.1582	-2.256		
+	0.1583	-2.194		
+	0.1584	-2.176		
+	0.1585	-2.144		
+	0.1586	-2.101		
+	0.1587	-1.933		
+	0.1588	-1.902		
+	0.1589	-2.014		
+	0.159	-1.84		
+	0.1591	-1.784		
+	0.1592	-1.809		
+	0.1593	-1.79		
+	0.1594	-1.703		
+	0.1595	-1.721		
+	0.1596	-1.759		
+	0.1597	-1.566		
+	0.1598	-1.491		
+	0.1599	-1.547		
+	0.16	-1.448		
+	0.1601	-1.361		
+	0.1602	-1.323		
+	0.1603	-1.149		
+	0.1604	-1		
+	0.1605	-1		
+	0.1606	-0.981		
+	0.1607	-0.813		
+	0.1608	-0.826		
+	0.1609	-0.844		
+	0.161	-0.708		
+	0.1611	-0.589		
+	0.1612	-0.664		
+	0.1613	-0.602		
+	0.1614	-0.44		
+	0.1615	-0.496		
+	0.1616	-0.54		
+	0.1617	-0.459		
+	0.1618	-0.403		
+	0.1619	-0.372		
+	0.162	-0.365		
+	0.1621	-0.197		
+	0.1622	-0.191		
+	0.1623	0.026		
+	0.1624	0.456		
+	0.1625	0.959		
+	0.1626	1.749		
+	0.1627	3.13		
+	0.1628	4.947		
+	0.1629	7.472		
+	0.163	10.545		
+	0.1631	14.122		
+	0.1632	17.798		
+	0.1633	21.965		
+	0.1634	26.637		
+	0.1635	31.433		
+	0.1636	36.558		
+	0.1637	42.169		
+	0.1638	48.109		
+	0.1639	54.037		
+	0.164	60.363		
+	0.1641	66.677		
+	0.1642	72.86		
+	0.1643	78.993		
+	0.1644	84.896		
+	0.1645	89.76		
+	0.1646	93.542		
+	0.1647	96.559		
+	0.1648	98.724		
+	0.1649	100.098		
+	0.165	101.168		
+	0.1651	102.039		
+	0.1652	102.537		
+	0.1653	103.016		
+	0.1654	103.675		
+	0.1655	104.253		
+	0.1656	104.851		
+	0.1657	105.653		
+	0.1658	106.555		
+	0.1659	107.189		
+	0.166	107.998		
+	0.1661	108.813		
+	0.1662	109.373		
+	0.1663	109.858		
+	0.1664	110.48		
+	0.1665	110.822		
+	0.1666	111.058		
+	0.1667	111.338		
+	0.1668	111.736		
+	0.1669	111.811		
+	0.167	112.029		
+	0.1671	112.278		
+	0.1672	112.259		
+	0.1673	112.246		
+	0.1674	112.489		
+	0.1675	112.526		
+	0.1676	112.414		
+	0.1677	112.545		
+	0.1678	112.595		
+	0.1679	112.477		
+	0.168	112.489		
+	0.1681	112.757		
+	0.1682	112.744		
+	0.1683	112.8		
+	0.1684	113.13		
+	0.1685	113.372		
+	0.1686	113.428		
+	0.1687	113.69		
+	0.1688	113.907		
+	0.1689	113.82		
+	0.169	113.714		
+	0.1691	113.547		
+	0.1692	113.005		
+	0.1693	112.159		
+	0.1694	110.872		
+	0.1695	108.962		
+	0.1696	106.175		
+	0.1697	102.742		
+	0.1698	97.716		
+	0.1699	89.853		
+	0.17	80.305		
+	0.1701	72.76		
+	0.1702	66.173		
+	0.1703	59.965		
+	0.1704	54.435		
+	0.1705	49.179		
+	0.1706	44.06		
+	0.1707	39.494		
+	0.1708	35.208		
+	0.1709	31.003		
+	0.171	27.259		
+	0.1711	23.701		
+	0.1712	20.292		
+	0.1713	17.064		
+	0.1714	14.364		
+	0.1715	11.714		
+	0.1716	9.189		
+	0.1717	7.043		
+	0.1718	5.27		
+	0.1719	3.497		
+	0.172	2.011		
+	0.1721	0.953		
+	0.1722	-0.104		
+	0.1723	-1.062		
+	0.1724	-1.566		
+	0.1725	-2.014		
+	0.1726	-2.449		
+	0.1727	-2.698		
+	0.1728	-2.804		
+	0.1729	-2.959		
+	0.173	-3.028		
+	0.1731	-2.922		
+	0.1732	-2.928		
+	0.1733	-2.984		
+	0.1734	-2.822		
+	0.1735	-2.704		
+	0.1736	-2.773		
+	0.1737	-2.623		
+	0.1738	-2.431		
+	0.1739	-2.487		
+	0.174	-2.462		
+	0.1741	-2.263		
+	0.1742	-2.238		
+	0.1743	-2.294		
+	0.1744	-2.163		
+	0.1745	-2.07		
+	0.1746	-2.176		
+	0.1747	-2.132		
+	0.1748	-2.02		
+	0.1749	-1.983		
+	0.175	-2.07		
+	0.1751	-1.958		
+	0.1752	-1.877		
+	0.1753	-1.933		
+	0.1754	-1.777		
+	0.1755	-1.659		
+	0.1756	-1.74		
+	0.1757	-1.665		
+	0.1758	-1.522		
+	0.1759	-1.572		
+	0.176	-1.547		
+	0.1761	-1.448		
+	0.1762	-1.398		
+	0.1763	-1.448		
+	0.1764	-1.28		
+	0.1765	-1.162		
+	0.1766	-1.274		
+	0.1767	-1.174		
+	0.1768	-0.981		
+	0.1769	-0.994		
+	0.177	-0.95		
+	0.1771	-0.714		
+	0.1772	-0.645		
+	0.1773	-0.695		
+	0.1774	-0.558		
+	0.1775	-0.459		
+	0.1776	-0.533		
+	0.1777	-0.509		
+	0.1778	-0.347		
+	0.1779	-0.403		
+	0.178	-0.502		
+	0.1781	-0.334		
+	0.1782	-0.347		
+	0.1783	-0.453		
+	0.1784	-0.303		
+	0.1785	-0.067		
+	0.1786	0.033		
+	0.1787	0.443		
+	0.1788	1.071		
+	0.1789	1.973		
+	0.179	3.255		
+	0.1791	5.301		
+	0.1792	8.032		
+	0.1793	10.974		
+	0.1794	14.408		
+	0.1795	18.37		
+	0.1796	22.469		
+	0.1797	26.998		
+	0.1798	31.968		
+	0.1799	37.155		
+	0.18	42.617		
+	0.1801	48.545		
+	0.1802	54.628		
+	0.1803	60.73		
+	0.1804	67.075		
+	0.1805	73.382		
+	0.1806	79.416		
+	0.1807	85.101		
+	0.1808	90.109		
+	0.1809	93.878		
+	0.181	96.64		
+	0.1811	98.773		
+	0.1812	100.297		
+	0.1813	101.243		
+	0.1814	101.983		
+	0.1815	102.649		
+	0.1816	103.04		
+	0.1817	103.463		
+	0.1818	104.229		
+	0.1819	104.869		
+	0.182	105.622		
+	0.1821	106.524		
+	0.1822	107.32		
+	0.1823	108.004		
+	0.1824	108.732		
+	0.1825	109.478		
+	0.1826	109.976		
+	0.1827	110.399		
+	0.1828	110.816		
+	0.1829	111.17		
+	0.183	111.332		
+	0.1831	111.687		
+	0.1832	111.898		
+	0.1833	111.879		
+	0.1834	112.147		
+	0.1835	112.296		
+	0.1836	112.321		
+	0.1837	112.358		
+	0.1838	112.564		
+	0.1839	112.557		
+	0.184	112.589		
+	0.1841	112.589		
+	0.1842	112.744		
+	0.1843	112.676		
+	0.1844	112.732		
+	0.1845	112.881		
+	0.1846	112.924		
+	0.1847	113.105		
+	0.1848	113.329		
+	0.1849	113.528		
+	0.185	113.584		
+	0.1851	113.77		
+	0.1852	113.851		
+	0.1853	113.814		
+	0.1854	113.515		
+	0.1855	113.136		
+	0.1856	112.253		
+	0.1857	110.915		
+	0.1858	109.18		
+	0.1859	106.592		
+	0.186	102.935		
+	0.1861	98.039		
+	0.1862	90.569		
+	0.1863	80.921		
+	0.1864	73.133		
+	0.1865	66.646		
+	0.1866	60.351		
+	0.1867	54.659		
+	0.1868	49.415		
+	0.1869	44.514		
+	0.187	39.836		
+	0.1871	35.463		
+	0.1872	31.507		
+	0.1873	27.62		
+	0.1874	23.943		
+	0.1875	20.734		
+	0.1876	17.599		
+	0.1877	14.601		
+	0.1878	11.988		
+	0.1879	9.537		
+	0.188	7.236		
+	0.1881	5.345		
+	0.1882	3.709		
+	0.1883	2.172		
+	0.1884	0.848		
+	0.1885	-0.054		
+	0.1886	-0.807		
+	0.1887	-1.572		
+	0.1888	-2.001		
+	0.1889	-2.343		
+	0.189	-2.636		
+	0.1891	-2.841		
+	0.1892	-2.81		
+	0.1893	-2.903		
+	0.1894	-2.966		
+	0.1895	-2.903		
+	0.1896	-2.847		
+	0.1897	-2.878		
+	0.1898	-2.816		
+	0.1899	-2.729		
+	0.19	-2.71		
+	0.1901	-2.667		
+	0.1902	-2.468		
+	0.1903	-2.418		
+	0.1904	-2.418		
+	0.1905	-2.263		
+	0.1906	-2.194		
+	0.1907	-2.2		
+	0.1908	-2.144		
+	0.1909	-2.001		
+	0.191	-2.045		
+	0.1911	-2.039		
+	0.1912	-1.952		
+	0.1913	-1.989		
+	0.1914	-2.008		
+	0.1915	-1.945		
+	0.1916	-1.877		
+	0.1917	-1.902		
+	0.1918	-1.827		
+	0.1919	-1.709		
+	0.192	-1.665		
+	0.1921	-1.609		
+	0.1922	-1.547		
+	0.1923	-1.466		
+	0.1924	-1.504		
+	0.1925	-1.323		
+	0.1926	-1.267		
+	0.1927	-1.249		
+	0.1928	-1.211		
+	0.1929	-1.099		
+	0.193	-1.131		
+	0.1931	-1.081		
+	0.1932	-0.956		
+	0.1933	-0.857		
+	0.1934	-0.851		
+	0.1935	-0.776		
+	0.1936	-0.602		
+	0.1937	-0.627		
+	0.1938	-0.453		
+	0.1939	-0.403		
+	0.194	-0.434		
+	0.1941	-0.403		
+	0.1942	-0.272		
+	0.1943	-0.297		
+	0.1944	-0.39		
+	0.1945	-0.272		
+	0.1946	-0.266		
+	0.1947	-0.272		
+	0.1948	-0.079		
+	0.1949	0.188		
+	0.195	0.536		
+	0.1951	1.165		
+	0.1952	2.235		
+	0.1953	3.715		
+	0.1954	5.836		
+	0.1955	8.778		
+	0.1956	11.907		
+	0.1957	15.403		
+	0.1958	19.316		
+	0.1959	23.738		
+	0.196	28.217		
+	0.1961	33.056		
+	0.1962	38.412		
+	0.1963	43.96		
+	0.1964	49.776		
+	0.1965	55.791		
+	0.1966	62.067		
+	0.1967	68.207		
+	0.1968	74.452		
+	0.1969	80.523		
+	0.197	86.14		
+	0.1971	90.687		
+	0.1972	94.313		
+	0.1973	97.025		
+	0.1974	98.948		
+	0.1975	100.384		
+	0.1976	101.355		
+	0.1977	102.027		
+	0.1978	102.562		
+	0.1979	103.028		
+	0.198	103.613		
+	0.1981	104.166		
+	0.1982	104.894		
+	0.1983	105.603		
+	0.1984	106.406		
+	0.1985	107.158		
+	0.1986	108.042		
+	0.1987	108.776		
+	0.1988	109.404		
+	0.1989	109.982		
+	0.199	110.461		
+	0.1991	110.735		
+	0.1992	111.251		
+	0.1993	111.457		
+	0.1994	111.662		
+	0.1995	111.724		
+	0.1996	111.942		
+	0.1997	112.072		
+	0.1998	112.041		
+	0.1999	112.222		
+	0.2	112.284		
+	0.2001	112.24		
+	0.2002	112.302		
+	0.2003	112.464		
+	0.2004	112.495		
+	0.2005	112.57		
+	0.2006	112.651		
+	0.2007	112.757		
+	0.2008	112.875		
+	0.2009	112.993		
+	0.201	113.161		
+	0.2011	113.323		
+	0.2012	113.422		
+	0.2013	113.665		
+	0.2014	113.708		
+	0.2015	113.64		
+	0.2016	113.596		
+	0.2017	113.329		
+	0.2018	112.701		
+	0.2019	111.923		
+	0.202	110.573		
+	0.2021	108.57		
+	0.2022	105.877		
+	0.2023	102.163		
+	0.2024	96.969		
+	0.2025	88.852		
+	0.2026	79.64		
+	0.2027	72.138		
+	0.2028	65.482		
+	0.2029	59.467		
+	0.203	53.944		
+	0.2031	48.681		
+	0.2032	43.687		
+	0.2033	39.146		
+	0.2034	34.848		
+	0.2035	30.823		
+	0.2036	27.103		
+	0.2037	23.589		
+	0.2038	20.224		
+	0.2039	17.163		
+	0.204	14.333		
+	0.2041	11.646		
+	0.2042	9.301		
+	0.2043	7.223		
+	0.2044	5.202		
+	0.2045	3.454		
+	0.2046	2.073		
+	0.2047	0.885		
+	0.2048	-0.173		
+	0.2049	-1.031		
+	0.205	-1.572		
+	0.2051	-2.107		
+	0.2052	-2.474		
+	0.2053	-2.605		
+	0.2054	-2.779		
+	0.2055	-2.86		
+	0.2056	-2.891		
+	0.2057	-2.86		
+	0.2058	-2.847		
+	0.2059	-2.829		
+	0.206	-2.692		
+	0.2061	-2.698		
+	0.2062	-2.704		
+	0.2063	-2.567		
+	0.2064	-2.611		
+	0.2065	-2.567		
+	0.2066	-2.412		
+	0.2067	-2.368		
+	0.2068	-2.387		
+	0.2069	-2.281		
+	0.207	-2.169		
+	0.2071	-2.113		
+	0.2072	-2.082		
+	0.2073	-1.989		
+	0.2074	-1.952		
+	0.2075	-1.976		
+	0.2076	-1.952		
+	0.2077	-1.84		
+	0.2078	-1.927		
+	0.2079	-1.858		
+	0.208	-1.809		
+	0.2081	-1.858		
+	0.2082	-1.846		
+	0.2083	-1.759		
+	0.2084	-1.653		
+	0.2085	-1.609		
+	0.2086	-1.504		
+	0.2087	-1.392		
+	0.2088	-1.386		
+	0.2089	-1.305		
+	0.209	-1.162		
+	0.2091	-1.131		
+	0.2092	-1.112		
+	0.2093	-0.981		
+	0.2094	-0.9		
+	0.2095	-0.975		
+	0.2096	-0.869		
+	0.2097	-0.751		
+	0.2098	-0.764		
+	0.2099	-0.72		
+	0.21	-0.54		
+	0.2101	-0.509		
+	0.2102	-0.533		
+	0.2103	-0.378		
+	0.2104	-0.291		
+	0.2105	-0.266		
+	0.2106	-0.26		
+	0.2107	-0.222		
+	0.2108	-0.26		
+	0.2109	-0.229		
+	0.211	-0.123		
+	0.2111	-0.042		
+	0.2112	0.039		
+	0.2113	0.53		
+	0.2114	1.215		
+	0.2115	1.961		
+	0.2116	3.429		
+	0.2117	5.674		
+	0.2118	8.331		
+	0.2119	11.497		
+	0.212	15.092		
+	0.2121	18.967		
+	0.2122	23.066		
+	0.2123	27.694		
+	0.2124	32.664		
+	0.2125	37.796		
+	0.2126	43.239		
+	0.2127	49.123		
+	0.2128	55.032		
+	0.2129	61.147		
+	0.213	67.448		
+	0.2131	73.637		
+	0.2132	79.546		
+	0.2133	85.232		
+	0.2134	90.021		
+	0.2135	93.642		
+	0.2136	96.497		
+	0.2137	98.587		
+	0.2138	100.073		
+	0.2139	101.044		
+	0.214	101.809		
+	0.2141	102.394		
+	0.2142	102.823		
+	0.2143	103.389		
+	0.2144	104.036		
+	0.2145	104.571		
+	0.2146	105.33		
+	0.2147	106.225		
+	0.2148	106.965		
+	0.2149	107.668		
+	0.215	108.433		
+	0.2151	109.13		
+	0.2152	109.615		
+	0.2153	110.113		
+	0.2154	110.691		
+	0.2155	110.984		
+	0.2156	111.195		
+	0.2157	111.556		
+	0.2158	111.718		
+	0.2159	111.724		
+	0.216	112.004		
+	0.2161	112.06		
+	0.2162	112.004		
+	0.2163	112.11		
+	0.2164	112.271		
+	0.2165	112.209		
+	0.2166	112.184		
+	0.2167	112.315		
+	0.2168	112.377		
+	0.2169	112.377		
+	0.217	112.551		
+	0.2171	112.769		
+	0.2172	112.806		
+	0.2173	112.962		
+	0.2174	113.229		
+	0.2175	113.36		
+	0.2176	113.441		
+	0.2177	113.634		
+	0.2178	113.615		
+	0.2179	113.416		
+	0.218	113.242		
+	0.2181	112.8		
+	0.2182	111.867		
+	0.2183	110.598		
+	0.2184	108.807		
+	0.2185	106.219		
+	0.2186	102.773		
+	0.2187	98.07		
+	0.2188	90.625		
+	0.2189	81.095		
+	0.219	73.42		
+	0.2191	66.913		
+	0.2192	60.674		
+	0.2193	54.995		
+	0.2194	49.807		
+	0.2195	44.707		
+	0.2196	39.936		
+	0.2197	35.781		
+	0.2198	31.688		
+	0.2199	27.713		
+	0.22	24.186		
+	0.2201	20.883		
+	0.2202	17.673		
+	0.2203	14.75		
+	0.2204	12.28		
+	0.2205	9.823		
+	0.2206	7.516		
+	0.2207	5.643		
+	0.2208	3.958		
+	0.2209	2.347		
+	0.221	1.165		
+	0.2211	0.089		
+	0.2212	-0.857		
+	0.2213	-1.572		
+	0.2214	-1.908		
+	0.2215	-2.399		
+	0.2216	-2.717		
+	0.2217	-2.773		
+	0.2218	-2.903		
+	0.2219	-2.959		
+	0.222	-2.847		
+	0.2221	-2.816		
+	0.2222	-2.872		
+	0.2223	-2.791		
+	0.2224	-2.611		
+	0.2225	-2.592		
+	0.2226	-2.673		
+	0.2227	-2.524		
+	0.2228	-2.474		
+	0.2229	-2.48		
+	0.223	-2.437		
+	0.2231	-2.337		
+	0.2232	-2.3		
+	0.2233	-2.281		
+	0.2234	-2.144		
+	0.2235	-2.144		
+	0.2236	-2.194		
+	0.2237	-1.958		
+	0.2238	-1.889		
+	0.2239	-1.976		
+	0.224	-1.939		
+	0.2241	-1.734		
+	0.2242	-1.802		
+	0.2243	-1.889		
+	0.2244	-1.709		
+	0.2245	-1.74		
+	0.2246	-1.821		
+	0.2247	-1.634		
+	0.2248	-1.541		
+	0.2249	-1.591		
+	0.225	-1.529		
+	0.2251	-1.404		
+	0.2252	-1.361		
+	0.2253	-1.342		
+	0.2254	-1.131		
+	0.2255	-0.981		
+	0.2256	-1.118		
+	0.2257	-0.919		
+	0.2258	-0.807		
+	0.2259	-0.832		
+	0.226	-0.739		
+	0.2261	-0.602		
+	0.2262	-0.614		
+	0.2263	-0.664		
+	0.2264	-0.477		
+	0.2265	-0.471		
+	0.2266	-0.583		
+	0.2267	-0.434		
+	0.2268	-0.409		
+	0.2269	-0.378		
+	0.227	-0.334		
+	0.2271	-0.135		
+	0.2272	-0.197		
+	0.2273	-0.266		
+	0.2274	0.014		
+	0.2275	0.306		
+	0.2276	0.555		
+	0.2277	1.302		
+	0.2278	2.303		
+	0.2279	3.609		
+	0.228	5.83		
+	0.2281	8.642		
+	0.2282	11.745		
+	0.2283	15.167		
+	0.2284	19.191		
+	0.2285	23.421		
+	0.2286	27.831		
+	0.2287	32.863		
+	0.2288	38.163		
+	0.2289	43.512		
+	0.229	49.31		
+	0.2291	55.374		
+	0.2292	61.439		
+	0.2293	67.485		
+	0.2294	73.637		
+	0.2295	79.646		
+	0.2296	85.139		
+	0.2297	89.909		
+	0.2298	93.654		
+	0.2299	96.279		
+	0.23	98.251		
+	0.2301	99.8		
+	0.2302	100.832		
+	0.2303	101.492		
+	0.2304	102.207		
+	0.2305	102.792		
+	0.2306	103.152		
+	0.2307	103.812		
+	0.2308	104.589		
+	0.2309	105.174		
+	0.231	105.976		
+	0.2311	106.841		
+	0.2312	107.625		
+	0.2313	108.166		
+	0.2314	108.9		
+	0.2315	109.547		
+	0.2316	109.883		
+	0.2317	110.505		
+	0.2318	110.735		
+	0.2319	110.971		
+	0.232	111.208		
+	0.2321	111.544		
+	0.2322	111.693		
+	0.2323	111.705		
+	0.2324	111.911		
+	0.2325	111.991		
+	0.2326	111.942		
+	0.2327	111.991		
+	0.2328	112.147		
+	0.2329	112.091		
+	0.233	112.066		
+	0.2331	112.246		
+	0.2332	112.184		
+	0.2333	112.191		
+	0.2334	112.701		
+	0.2335	112.663		
+	0.2336	112.669		
+	0.2337	112.9		
+	0.2338	113.198		
+	0.2339	113.291		
+	0.234	113.279		
+	0.2341	113.459		
+	0.2342	113.347		
+	0.2343	113.03		
+	0.2344	112.495		
+	0.2345	111.68		
+	0.2346	110.287		
+	0.2347	108.44		
+	0.2348	105.964		
+	0.2349	102.356		
+	0.235	97.361		
+	0.2351	89.878		
+	0.2352	80.647		
+	0.2353	72.841		
+	0.2354	66.428		
+	0.2355	60.419		
+	0.2356	54.703		
+	0.2357	49.409		
+	0.2358	44.676		
+	0.2359	39.892		
+	0.236	35.482		
+	0.2361	31.538		
+	0.2362	27.719		
+	0.2363	23.975		
+	0.2364	20.721		
+	0.2365	17.698		
+	0.2366	14.657		
+	0.2367	11.982		
+	0.2368	9.668		
+	0.2369	7.491		
+	0.237	5.494		
+	0.2371	3.877		
+	0.2372	2.434		
+	0.2373	1.047		
+	0.2374	0.064		
+	0.2375	-0.695		
+	0.2376	-1.466		
+	0.2377	-2.02		
+	0.2378	-2.312		
+	0.2379	-2.636		
+	0.238	-2.928		
+	0.2381	-2.841		
+	0.2382	-2.891		
+	0.2383	-2.99		
+	0.2384	-2.953		
+	0.2385	-2.829		
+	0.2386	-2.847		
+	0.2387	-2.729		
+	0.2388	-2.543		
+	0.2389	-2.586		
+	0.239	-2.524		
+	0.2391	-2.424		
+	0.2392	-2.35		
+	0.2393	-2.356		
+	0.2394	-2.356		
+	0.2395	-2.25		
+	0.2396	-2.306		
+	0.2397	-2.219		
+	0.2398	-2.138		
+	0.2399	-2.088		
+	0.24	-2.101		
+	0.2401	-2.045		
+	0.2402	-1.896		
+	0.2403	-1.939		
+	0.2404	-1.852		
+	0.2405	-1.79		
+	0.2406	-1.802		
+	0.2407	-1.846		
+	0.2408	-1.609		
+	0.2409	-1.653		
+	0.241	-1.672		
+	0.2411	-1.634		
+	0.2412	-1.554		
+	0.2413	-1.578		
+	0.2414	-1.442		
+	0.2415	-1.311		
+	0.2416	-1.342		
+	0.2417	-1.348		
+	0.2418	-1.149		
+	0.2419	-1.025		
+	0.242	-1.006		
+	0.2421	-0.844		
+	0.2422	-0.77		
+	0.2423	-0.751		
+	0.2424	-0.664		
+	0.2425	-0.459		
+	0.2426	-0.502		
+	0.2427	-0.527		
+	0.2428	-0.409		
+	0.2429	-0.428		
+	0.243	-0.459		
+	0.2431	-0.397		
+	0.2432	-0.328		
+	0.2433	-0.365		
+	0.2434	-0.372		
+	0.2435	-0.173		
+	0.2436	-0.185		
+	0.2437	-0.067		
+	0.2438	0.194		
+	0.2439	0.574		
+	0.244	1.115		
+	0.2441	2.073		
+	0.2442	3.528		
+	0.2443	5.556		
+	0.2444	8.144		
+	0.2445	11.291		
+	0.2446	14.632		
+	0.2447	18.37		
+	0.2448	22.618		
+	0.2449	27.134		
+	0.245	31.837		
+	0.2451	37.018		
+	0.2452	42.511		
+	0.2453	48.234		
+	0.2454	54.099		
+	0.2455	60.332		
+	0.2456	66.328		
+	0.2457	72.343		
+	0.2458	78.421		
+	0.2459	84.087		
+	0.246	88.883		
+	0.2461	92.733		
+	0.2462	95.657		
+	0.2463	97.716		
+	0.2464	99.29		
+	0.2465	100.447		
+	0.2466	101.224		
+	0.2467	101.734		
+	0.2468	102.375		
+	0.2469	102.966		
+	0.247	103.463		
+	0.2471	104.173		
+	0.2472	104.919		
+	0.2473	105.74		
+	0.2474	106.487		
+	0.2475	107.376		
+	0.2476	108.085		
+	0.2477	108.626		
+	0.2478	109.205		
+	0.2479	109.74		
+	0.248	110.082		
+	0.2481	110.492		
+	0.2482	110.81		
+	0.2483	111.009		
+	0.2484	111.139		
+	0.2485	111.394		
+	0.2486	111.562		
+	0.2487	111.693		
+	0.2488	111.774		
+	0.2489	111.879		
+	0.249	111.96		
+	0.2491	111.929		
+	0.2492	112.041		
+	0.2493	112.06		
+	0.2494	111.985		
+	0.2495	112.091		
+	0.2496	112.103		
+	0.2497	112.228		
+	0.2498	112.358		
+	0.2499	112.595		
+	0.25	112.669		
+	0.2501	112.837		
+	0.2502	113.03		
+	0.2503	113.242		
+	0.2504	113.211		
+	0.2505	113.167		
+	0.2506	113.018		
+	0.2507	112.539		
+	0.2508	111.824		
+	0.2509	110.673		
+	0.251	108.863		
+	0.2511	106.449		
+	0.2512	103.296		
+	0.2513	98.599		
+	0.2514	91.85		
+	0.2515	82.551		
+	0.2516	74.458		
+	0.2517	67.628		
+	0.2518	61.62		
+	0.2519	55.959		
+	0.252	50.697		
+	0.2521	45.665		
+	0.2522	40.925		
+	0.2523	36.62		
+	0.2524	32.484		
+	0.2525	28.59		
+	0.2526	25.063		
+	0.2527	21.598		
+	0.2528	18.37		
+	0.2529	15.496		
+	0.253	12.691		
+	0.2531	10.215		
+	0.2532	8.044		
+	0.2533	5.998		
+	0.2534	4.2		
+	0.2535	2.639		
+	0.2536	1.42		
+	0.2537	0.356		
+	0.2538	-0.577		
+	0.2539	-1.236		
+	0.254	-1.765		
+	0.2541	-2.232		
+	0.2542	-2.399		
+	0.2543	-2.673		
+	0.2544	-2.81		
+	0.2545	-2.928		
+	0.2546	-2.903		
+	0.2547	-2.86		
+	0.2548	-2.922		
+	0.2549	-2.76		
+	0.255	-2.773		
+	0.2551	-2.748		
+	0.2552	-2.667		
+	0.2553	-2.449		
+	0.2554	-2.455		
+	0.2555	-2.381		
+	0.2556	-2.306		
+	0.2557	-2.25		
+	0.2558	-2.219		
+	0.2559	-2.169		
+	0.256	-2.101		
+	0.2561	-2.107		
+	0.2562	-2.101		
+	0.2563	-2.07		
+	0.2564	-2.032		
+	0.2565	-2.008		
+	0.2566	-1.939		
+	0.2567	-1.989		
+	0.2568	-1.952		
+	0.2569	-1.79		
+	0.257	-1.709		
+	0.2571	-1.715		
+	0.2572	-1.672		
+	0.2573	-1.522		
+	0.2574	-1.547		
+	0.2575	-1.529		
+	0.2576	-1.392		
+	0.2577	-1.392		
+	0.2578	-1.379		
+	0.2579	-1.255		
+	0.258	-1.224		
+	0.2581	-1.168		
+	0.2582	-1.081		
+	0.2583	-1.012		
+	0.2584	-0.913		
+	0.2585	-0.888		
+	0.2586	-0.726		
+	0.2587	-0.627		
+	0.2588	-0.558		
+	0.2589	-0.44		
+	0.259	-0.365		
+	0.2591	-0.397		
+	0.2592	-0.229		
+	0.2593	-0.185		
+	0.2594	-0.21		
+	0.2595	-0.322		
+	0.2596	-0.316		
+	0.2597	-0.241		
+	0.2598	-0.278		
+	0.2599	-0.123		
+	0.26	-0.16		
+	0.2601	0.07		
+	0.2602	0.344		
+	0.2603	1.003		
+	0.2604	1.743		
+	0.2605	3.068		
+	0.2606	4.828		
+	0.2607	7.397		
+	0.2608	10.277		
+	0.2609	13.593		
+	0.261	17.306		
+	0.2611	21.3		
+	0.2612	25.66		
+	0.2613	30.276		
+	0.2614	35.271		
+	0.2615	40.539		
+	0.2616	46.137		
+	0.2617	51.972		
+	0.2618	57.999		
+	0.2619	64.07		
+	0.262	70.26		
+	0.2621	76.212		
+	0.2622	81.96		
+	0.2623	87.185		
+	0.2624	91.409		
+	0.2625	94.606		
+	0.2626	97.044		
+	0.2627	98.748		
+	0.2628	99.993		
+	0.2629	100.832		
+	0.263	101.517		
+	0.2631	102.045		
+	0.2632	102.512		
+	0.2633	103.208		
+	0.2634	103.774		
+	0.2635	104.44		
+	0.2636	105.305		
+	0.2637	106.175		
+	0.2638	106.959		
+	0.2639	107.662		
+	0.264	108.39		
+	0.2641	108.999		
+	0.2642	109.609		
+	0.2643	110.057		
+	0.2644	110.38		
+	0.2645	110.617		
+	0.2646	110.928		
+	0.2647	111.214		
+	0.2648	111.301		
+	0.2649	111.481		
+	0.265	111.562		
+	0.2651	111.643		
+	0.2652	111.662		
+	0.2653	111.892		
+	0.2654	111.935		
+	0.2655	111.873		
+	0.2656	111.998		
+	0.2657	112.091		
+	0.2658	112.079		
+	0.2659	112.141		
+	0.266	112.271		
+	0.2661	112.383		
+	0.2662	112.408		
+	0.2663	112.645		
+	0.2664	112.831		
+	0.2665	112.949		
+	0.2666	113.092		
+	0.2667	113.167		
+	0.2668	113.148		
+	0.2669	113.018		
+	0.267	112.757		
+	0.2671	112.166		
+	0.2672	111.096		
+	0.2673	109.628		
+	0.2674	107.569		
+	0.2675	104.571		
+	0.2676	100.621		
+	0.2677	95.041		
+	0.2678	86.215		
+	0.2679	77.369		
+	0.268	70.372		
+	0.2681	64.126		
+	0.2682	58.149		
+	0.2683	52.718		
+	0.2684	47.699		
+	0.2685	42.729		
+	0.2686	38.374		
+	0.2687	34.244		
+	0.2688	30.232		
+	0.2689	26.531		
+	0.269	23.023		
+	0.2691	19.801		
+	0.2692	16.778		
+	0.2693	13.985		
+	0.2694	11.403		
+	0.2695	8.946		
+	0.2696	6.875		
+	0.2697	5.04		
+	0.2698	3.379		
+	0.2699	1.861		
+	0.27	0.76		
+	0.2701	-0.222		
+	0.2702	-1.099		
+	0.2703	-1.578		
+	0.2704	-1.989		
+	0.2705	-2.319		
+	0.2706	-2.605		
+	0.2707	-2.648		
+	0.2708	-2.723		
+	0.2709	-2.86		
+	0.271	-2.785		
+	0.2711	-2.723		
+	0.2712	-2.829		
+	0.2713	-2.773		
+	0.2714	-2.623		
+	0.2715	-2.679		
+	0.2716	-2.679		
+	0.2717	-2.511		
+	0.2718	-2.505		
+	0.2719	-2.449		
+	0.272	-2.275		
+	0.2721	-2.157		
+	0.2722	-2.275		
+	0.2723	-2.138		
+	0.2724	-2.045		
+	0.2725	-2.008		
+	0.2726	-2.001		
+	0.2727	-1.896		
+	0.2728	-1.952		
+	0.2729	-1.958		
+	0.273	-1.858		
+	0.2731	-1.846		
+	0.2732	-1.883		
+	0.2733	-1.896		
+	0.2734	-1.709		
+	0.2735	-1.753		
+	0.2736	-1.684		
+	0.2737	-1.522		
+	0.2738	-1.435		
+	0.2739	-1.541		
+	0.274	-1.317		
+	0.2741	-1.187		
+	0.2742	-1.249		
+	0.2743	-1.23		
+	0.2744	-1.037		
+	0.2745	-1.081		
+	0.2746	-1.05		
+	0.2747	-0.9		
+	0.2748	-0.813		
+	0.2749	-0.882		
+	0.275	-0.714		
+	0.2751	-0.664		
+	0.2752	-0.639		
+	0.2753	-0.49		
+	0.2754	-0.353		
+	0.2755	-0.297		
+	0.2756	-0.365		
+	0.2757	-0.235		
+	0.2758	-0.173		
+	0.2759	-0.179		
+	0.276	-0.191		
+	0.2761	-0.098		
+	0.2762	-0.266		
+	0.2763	-0.166		
+	0.2764	0.101		
+	0.2765	0.263		
+	0.2766	0.624		
+	0.2767	1.382		
+	0.2768	2.471		
+	0.2769	4.001		
+	0.277	6.352		
+	0.2771	9.195		
+	0.2772	12.243		
+	0.2773	15.776		
+	0.2774	19.832		
+	0.2775	24.024		
+	0.2776	28.385		
+	0.2777	33.348		
+	0.2778	38.511		
+	0.2779	43.805		
+	0.278	49.621		
+	0.2781	55.592		
+	0.2782	61.526		
+	0.2783	67.492		
+	0.2784	73.569		
+	0.2785	79.422		
+	0.2786	84.883		
+	0.2787	89.592		
+	0.2788	93.312		
+	0.2789	95.831		
+	0.279	98.039		
+	0.2791	99.514		
+	0.2792	100.49		
+	0.2793	101.187		
+	0.2794	101.877		
+	0.2795	102.319		
+	0.2796	102.798		
+	0.2797	103.482		
+	0.2798	104.173		
+	0.2799	104.819		
+	0.28	105.578		
+	0.2801	106.487		
+	0.2802	107.283		
+	0.2803	107.973		
+	0.2804	108.8		
+	0.2805	109.366		
+	0.2806	109.69		
+	0.2807	110.206		
+	0.2808	110.617		
+	0.2809	110.778		
+	0.281	111.09		
+	0.2811	111.295		
+	0.2812	111.313		
+	0.2813	111.413		
+	0.2814	111.631		
+	0.2815	111.674		
+	0.2816	111.687		
+	0.2817	111.755		
+	0.2818	111.855		
+	0.2819	111.886		
+	0.282	111.948		
+	0.2821	112.228		
+	0.2822	112.122		
+	0.2823	112.116		
+	0.2824	112.377		
+	0.2825	112.464		
+	0.2826	112.483		
+	0.2827	112.744		
+	0.2828	113.012		
+	0.2829	112.993		
+	0.283	113.099		
+	0.2831	113.304		
+	0.2832	113.005		
+	0.2833	112.75		
+	0.2834	112.365		
+	0.2835	111.587		
+	0.2836	110.287		
+	0.2837	108.539		
+	0.2838	106.126		
+	0.2839	102.611		
+	0.284	97.89		
+	0.2841	90.799		
+	0.2842	81.425		
+	0.2843	73.581		
+	0.2844	67.125		
+	0.2845	61.085		
+	0.2846	55.331		
+	0.2847	50.087		
+	0.2848	45.223		
+	0.2849	40.452		
+	0.285	36.079		
+	0.2851	32.204		
+	0.2852	28.391		
+	0.2853	24.764		
+	0.2854	21.505		
+	0.2855	18.358		
+	0.2856	15.297		
+	0.2857	12.672		
+	0.2858	10.246		
+	0.2859	7.976		
+	0.286	5.948		
+	0.2861	4.262		
+	0.2862	2.627		
+	0.2863	1.239		
+	0.2864	0.325		
+	0.2865	-0.583		
+	0.2866	-1.423		
+	0.2867	-1.933		
+	0.2868	-2.244		
+	0.2869	-2.511		
+	0.287	-2.735		
+	0.2871	-2.679		
+	0.2872	-2.804		
+	0.2873	-2.835		
+	0.2874	-2.791		
+	0.2875	-2.611		
+	0.2876	-2.76		
+	0.2877	-2.661		
+	0.2878	-2.493		
+	0.2879	-2.623		
+	0.288	-2.642		
+	0.2881	-2.449		
+	0.2882	-2.406		
+	0.2883	-2.443		
+	0.2884	-2.281		
+	0.2885	-2.25		
+	0.2886	-2.194		
+	0.2887	-2.188		
+	0.2888	-1.933		
+	0.2889	-1.983		
+	0.289	-1.97		
+	0.2891	-1.771		
+	0.2892	-1.777		
+	0.2893	-1.889		
+	0.2894	-1.84		
+	0.2895	-1.777		
+	0.2896	-1.902		
+	0.2897	-1.796		
+	0.2898	-1.665		
+	0.2899	-1.678		
+	0.29	-1.753		
+	0.2901	-1.522		
+	0.2902	-1.417		
+	0.2903	-1.46		
+	0.2904	-1.249		
+	0.2905	-1.193		
+	0.2906	-1.211		
+	0.2907	-1.155		
+	0.2908	-0.925		
+	0.2909	-0.944		
+	0.291	-0.919		
+	0.2911	-0.857		
+	0.2912	-0.82		
+	0.2913	-0.757		
+	0.2914	-0.714		
+	0.2915	-0.552		
+	0.2916	-0.54		
+	0.2917	-0.577		
+	0.2918	-0.353		
+	0.2919	-0.285		
+	0.292	-0.334		
+	0.2921	-0.129		
+	0.2922	-0.191		
+	0.2923	-0.166		
+	0.2924	-0.123		
+	0.2925	-0.061		
+	0.2926	-0.03		
+	0.2927	-0.017		
+	0.2928	0.281		
+	0.2929	0.487		
+	0.293	1.04		
+	0.2931	2.017		
+	0.2932	3.385		
+	0.2933	5.258		
+	0.2934	8.032		
+	0.2935	11.061		
+	0.2936	14.364		
+	0.2937	18.127		
+	0.2938	22.401		
+	0.2939	26.668		
+	0.294	31.333		
+	0.2941	36.428		
+	0.2942	41.802		
+	0.2943	47.282		
+	0.2944	53.092		
+	0.2945	59.044		
+	0.2946	64.979		
+	0.2947	70.962		
+	0.2948	76.915		
+	0.2949	82.495		
+	0.295	87.477		
+	0.2951	91.676		
+	0.2952	94.823		
+	0.2953	96.945		
+	0.2954	98.761		
+	0.2955	100.16		
+	0.2956	100.894		
+	0.2957	101.56		
+	0.2958	102.188		
+	0.2959	102.611		
+	0.296	103.152		
+	0.2961	103.806		
+	0.2962	104.508		
+	0.2963	105.162		
+	0.2964	106.02		
+	0.2965	106.897		
+	0.2966	107.55		
+	0.2967	108.16		
+	0.2968	108.981		
+	0.2969	109.553		
+	0.297	109.933		
+	0.2971	110.405		
+	0.2972	110.729		
+	0.2973	110.866		
+	0.2974	111.17		
+	0.2975	111.469		
+	0.2976	111.525		
+	0.2977	111.593		
+	0.2978	111.724		
+	0.2979	111.78		
+	0.298	111.712		
+	0.2981	111.867		
+	0.2982	111.904		
+	0.2983	111.836		
+	0.2984	111.892		
+	0.2985	112.147		
+	0.2986	112.172		
+	0.2987	112.234		
+	0.2988	112.52		
+	0.2989	112.595		
+	0.299	112.676		
+	0.2991	112.974		
+	0.2992	113.186		
+	0.2993	113.242		
+	0.2994	113.18		
+	0.2995	113.242		
+	0.2996	113.024		
+	0.2997	112.582		
+	0.2998	111.991		
+	0.2999	110.94		
+	0.3	109.279		
+	0.3001	107.245		
+	0.3002	104.428		
+	0.3003	100.285		
+	0.3004	94.668		
+	0.3005	85.953		
+	0.3006	77.282		
+	0.3007	70.297		
+	0.3008	64.083		
+	0.3009	58.298		
+	0.301	52.824		
+	0.3011	47.724		
+	0.3012	43.002		
+	0.3013	38.374		
+	0.3014	34.232		
+	0.3015	30.332		
+	0.3016	26.562		
+	0.3017	23.004		
+	0.3018	19.913		
+	0.3019	16.902		
+	0.302	14.041		
+	0.3021	11.528		
+	0.3022	9.27		
+	0.3023	7.062		
+	0.3024	5.177		
+	0.3025	3.628		
+	0.3026	2.135		
+	0.3027	0.854		
+	0.3028	-0.104		
+	0.3029	-0.9		
+	0.303	-1.659		
+	0.3031	-2.076		
+	0.3032	-2.3		
+	0.3033	-2.686		
+	0.3034	-2.866		
+	0.3035	-2.847		
+	0.3036	-2.86		
+	0.3037	-2.86		
+	0.3038	-2.773		
+	0.3039	-2.673		
+	0.304	-2.679		
+	0.3041	-2.648		
+	0.3042	-2.511		
+	0.3043	-2.549		
+	0.3044	-2.543		
+	0.3045	-2.418		
+	0.3046	-2.325		
+	0.3047	-2.343		
+	0.3048	-2.281		
+	0.3049	-2.263		
+	0.305	-2.256		
+	0.3051	-2.238		
+	0.3052	-2.051		
+	0.3053	-1.976		
+	0.3054	-1.945		
+	0.3055	-1.796		
+	0.3056	-1.784		
+	0.3057	-1.821		
+	0.3058	-1.74		
+	0.3059	-1.709		
+	0.306	-1.784		
+	0.3061	-1.746		
+	0.3062	-1.628		
+	0.3063	-1.703		
+	0.3064	-1.659		
+	0.3065	-1.504		
+	0.3066	-1.417		
+	0.3067	-1.491		
+	0.3068	-1.373		
+	0.3069	-1.249		
+	0.307	-1.211		
+	0.3071	-1.062		
+	0.3072	-0.931		
+	0.3073	-0.801		
+	0.3074	-0.782		
+	0.3075	-0.652		
+	0.3076	-0.571		
+	0.3077	-0.596		
+	0.3078	-0.577		
+	0.3079	-0.471		
+	0.308	-0.477		
+	0.3081	-0.465		
+	0.3082	-0.353		
+	0.3083	-0.285		
+	0.3084	-0.403		
+	0.3085	-0.154		
+	0.3086	-0.179		
+	0.3087	-0.129		
+	0.3088	-0.104		
+	0.3089	0.008		
+	0.309	0.051		
+	0.3091	0.163		
+	0.3092	0.574		
+	0.3093	0.922		
+	0.3094	1.588		
+	0.3095	2.745		
+	0.3096	4.449		
+	0.3097	6.813		
+	0.3098	9.649		
+	0.3099	12.853		
+	0.31	16.404		
+	0.3101	20.298		
+	0.3102	24.696		
+	0.3103	29.224		
+	0.3104	34.089		
+	0.3105	39.264		
+	0.3106	44.775		
+	0.3107	50.423		
+	0.3108	56.289		
+	0.3109	62.217		
+	0.311	68.182		
+	0.3111	73.998		
+	0.3112	79.851		
+	0.3113	85.194		
+	0.3114	89.686		
+	0.3115	93.25		
+	0.3116	95.949		
+	0.3117	97.865		
+	0.3118	99.339		
+	0.3119	100.503		
+	0.312	101.286		
+	0.3121	101.865		
+	0.3122	102.45		
+	0.3123	103.016		
+	0.3124	103.501		
+	0.3125	104.21		
+	0.3126	104.994		
+	0.3127	105.678		
+	0.3128	106.362		
+	0.3129	107.239		
+	0.313	107.905		
+	0.3131	108.57		
+	0.3132	109.242		
+	0.3133	109.709		
+	0.3134	110.125		
+	0.3135	110.511		
+	0.3136	110.853		
+	0.3137	111.083		
+	0.3138	111.357		
+	0.3139	111.525		
+	0.314	111.575		
+	0.3141	111.724		
+	0.3142	111.879		
+	0.3143	111.96		
+	0.3144	111.879		
+	0.3145	111.848		
+	0.3146	111.991		
+	0.3147	112.035		
+	0.3148	111.985		
+	0.3149	112.11		
+	0.315	112.228		
+	0.3151	112.215		
+	0.3152	112.483		
+	0.3153	112.676		
+	0.3154	112.918		
+	0.3155	113.068		
+	0.3156	113.273		
+	0.3157	113.385		
+	0.3158	113.267		
+	0.3159	113.304		
+	0.316	113.117		
+	0.3161	112.452		
+	0.3162	111.68		
+	0.3163	110.461		
+	0.3164	108.62		
+	0.3165	106.138		
+	0.3166	102.779		
+	0.3167	98.058		
+	0.3168	91.066		
+	0.3169	81.904		
+	0.317	74.166		
+	0.3171	67.666		
+	0.3172	61.632		
+	0.3173	56.052		
+	0.3174	50.803		
+	0.3175	45.864		
+	0.3176	41.211		
+	0.3177	36.782		
+	0.3178	32.689		
+	0.3179	28.913		
+	0.318	25.331		
+	0.3181	21.86		
+	0.3182	18.681		
+	0.3183	15.789		
+	0.3184	13.052		
+	0.3185	10.557		
+	0.3186	8.343		
+	0.3187	6.346		
+	0.3188	4.567		
+	0.3189	2.981		
+	0.319	1.718		
+	0.3191	0.518		
+	0.3192	-0.378		
+	0.3193	-1.056		
+	0.3194	-1.765		
+	0.3195	-2.2		
+	0.3196	-2.505		
+	0.3197	-2.592		
+	0.3198	-2.847		
+	0.3199	-2.916		
+	0.32	-2.854		
+	0.3201	-2.841		
+	0.3202	-2.779		
+	0.3203	-2.667		
+	0.3204	-2.642		
+	0.3205	-2.555		
+	0.3206	-2.561		
+	0.3207	-2.356		
+	0.3208	-2.431		
+	0.3209	-2.381		
+	0.321	-2.238		
+	0.3211	-2.232		
+	0.3212	-2.281		
+	0.3213	-2.219		
+	0.3214	-2.113		
+	0.3215	-2.113		
+	0.3216	-2.101		
+	0.3217	-2.039		
+	0.3218	-1.989		
+	0.3219	-1.933		
+	0.322	-1.777		
+	0.3221	-1.759		
+	0.3222	-1.802		
+	0.3223	-1.634		
+	0.3224	-1.597		
+	0.3225	-1.622		
+	0.3226	-1.479		
+	0.3227	-1.491		
+	0.3228	-1.498		
+	0.3229	-1.473		
+	0.323	-1.448		
+	0.3231	-1.404		
+	0.3232	-1.361		
+	0.3233	-1.267		
+	0.3234	-1.062		
+	0.3235	-1.068		
+	0.3236	-0.938		
+	0.3237	-0.788		
+	0.3238	-0.708		
+	0.3239	-0.739		
+	0.324	-0.509		
+	0.3241	-0.49		
+	0.3242	-0.415		
+	0.3243	-0.278		
+	0.3244	-0.297		
+	0.3245	-0.322		
+	0.3246	-0.303		
+	0.3247	-0.222		
+	0.3248	-0.222		
+	0.3249	-0.235		
+	0.325	-0.179		
+	0.3251	-0.067		
+	0.3252	-0.216		
+	0.3253	0.039		
+	0.3254	0.219		
+	0.3255	0.344		
+	0.3256	0.717		
+	0.3257	1.382		
+	0.3258	2.222		
+	0.3259	3.678		
+	0.326	5.768		
+	0.3261	8.399		
+	0.3262	11.366		
+	0.3263	14.688		
+	0.3264	18.557		
+	0.3265	22.563		
+	0.3266	26.904		
+	0.3267	31.588		
+	0.3268	36.726		
+	0.3269	41.939		
+	0.327	47.636		
+	0.3271	53.421		
+	0.3272	59.212		
+	0.3273	65.184		
+	0.3274	71.249		
+	0.3275	76.99		
+	0.3276	82.576		
+	0.3277	87.533		
+	0.3278	91.595		
+	0.3279	94.568		
+	0.328	96.87		
+	0.3281	98.736		
+	0.3282	99.862		
+	0.3283	100.857		
+	0.3284	101.51		
+	0.3285	102.095		
+	0.3286	102.58		
+	0.3287	103.302		
+	0.3288	103.862		
+	0.3289	104.527		
+	0.329	105.386		
+	0.3291	106.2		
+	0.3292	106.872		
+	0.3293	107.693		
+	0.3294	108.396		
+	0.3295	108.968		
+	0.3296	109.454		
+	0.3297	110.076		
+	0.3298	110.393		
+	0.3299	110.635		
+	0.33	111.015		
+	0.3301	111.251		
+	0.3302	111.388		
+	0.3303	111.668		
+	0.3304	111.848		
+	0.3305	111.892		
+	0.3306	111.917		
+	0.3307	112.122		
+	0.3308	112.11		
+	0.3309	112.085		
+	0.331	112.24		
+	0.3311	112.215		
+	0.3312	112.153		
+	0.3313	112.203		
+	0.3314	112.402		
+	0.3315	112.514		
+	0.3316	112.607		
+	0.3317	112.837		
+	0.3318	113.074		
+	0.3319	113.18		
+	0.332	113.447		
+	0.3321	113.553		
+	0.3322	113.478		
+	0.3323	113.323		
+	0.3324	113.099		
+	0.3325	112.427		
+	0.3326	111.438		
+	0.3327	109.951		
+	0.3328	107.886		
+	0.3329	104.994		
+	0.333	101.199		
+	0.3331	95.993		
+	0.3332	87.508		
+	0.3333	78.701		
+	0.3334	71.703		
+	0.3335	65.433		
+	0.3336	59.443		
+	0.3337	54.186		
+	0.3338	49.117		
+	0.3339	44.147		
+	0.334	39.724		
+	0.3341	35.575		
+	0.3342	31.513		
+	0.3343	27.738		
+	0.3344	24.254		
+	0.3345	20.883		
+	0.3346	17.642		
+	0.3347	14.936		
+	0.3348	12.293		
+	0.3349	9.718		
+	0.335	7.609		
+	0.3351	5.755		
+	0.3352	3.951		
+	0.3353	2.477		
+	0.3354	1.407		
+	0.3355	0.281		
+	0.3356	-0.596		
+	0.3357	-1.143		
+	0.3358	-1.672		
+	0.3359	-2.207		
+	0.336	-2.406		
+	0.3361	-2.605		
+	0.3362	-2.816		
+	0.3363	-2.891		
+	0.3364	-2.754		
+	0.3365	-2.791		
+	0.3366	-2.866		
+	0.3367	-2.766		
+	0.3368	-2.611		
+	0.3369	-2.63		
+	0.337	-2.443		
+	0.3371	-2.35		
+	0.3372	-2.343		
+	0.3373	-2.269		
+	0.3374	-2.188		
+	0.3375	-2.138		
+	0.3376	-2.157		
+	0.3377	-2.088		
+	0.3378	-2.045		
+	0.3379	-2.057		
+	0.338	-2.07		
+	0.3381	-1.871		
+	0.3382	-1.914		
+	0.3383	-1.952		
+	0.3384	-1.79		
+	0.3385	-1.771		
+	0.3386	-1.883		
+	0.3387	-1.634		
+	0.3388	-1.498		
+	0.3389	-1.554		
+	0.339	-1.547		
+	0.3391	-1.33		
+	0.3392	-1.305		
+	0.3393	-1.342		
+	0.3394	-1.218		
+	0.3395	-1.211		
+	0.3396	-1.305		
+	0.3397	-1.068		
+	0.3398	-1.043		
+	0.3399	-1.012		
+	0.34	-0.956		
+	0.3401	-0.739		
+	0.3402	-0.67		
+	0.3403	-0.664		
+	0.3404	-0.397		
+	0.3405	-0.347		
+	0.3406	-0.39		
+	0.3407	-0.278		
+	0.3408	-0.104		
+	0.3409	-0.229		
+	0.341	-0.197		
+	0.3411	-0.067		
+	0.3412	-0.16		
+	0.3413	-0.26		
+	0.3414	-0.023		
+	0.3415	-0.017		
+	0.3416	-0.16		
+	0.3417	-0.104		
+	0.3418	0.25		
+	0.3419	0.418		
+	0.342	0.922		
+	0.3421	1.855		
+	0.3422	2.813		
+	0.3423	4.468		
+	0.3424	6.881		
+	0.3425	9.736		
+	0.3426	12.797		
+	0.3427	16.286		
+	0.3428	20.28		
+	0.3429	24.366		
+	0.343	28.764		
+	0.3431	33.678		
+	0.3432	38.692		
+	0.3433	44.035		
+	0.3434	49.801		
+	0.3435	55.648		
+	0.3436	61.433		
+	0.3437	67.479		
+	0.3438	73.463		
+	0.3439	79.08		
+	0.344	84.46		
+	0.3441	89.275		
+	0.3442	92.945		
+	0.3443	95.576		
+	0.3444	97.766		
+	0.3445	99.296		
+	0.3446	100.285		
+	0.3447	101.174		
+	0.3448	101.933		
+	0.3449	102.294		
+	0.345	102.736		
+	0.3451	103.526		
+	0.3452	104.123		
+	0.3453	104.77		
+	0.3454	105.703		
+	0.3455	106.53		
+	0.3456	107.177		
+	0.3457	108.004		
+	0.3458	108.701		
+	0.3459	109.261		
+	0.346	109.709		
+	0.3461	110.3		
+	0.3462	110.673		
+	0.3463	110.853		
+	0.3464	111.27		
+	0.3465	111.525		
+	0.3466	111.587		
+	0.3467	111.68		
+	0.3468	111.929		
+	0.3469	111.948		
+	0.347	112.06		
+	0.3471	112.228		
+	0.3472	112.253		
+	0.3473	112.166		
+	0.3474	112.321		
+	0.3475	112.495		
+	0.3476	112.464		
+	0.3477	112.508		
+	0.3478	112.682		
+	0.3479	112.738		
+	0.348	112.844		
+	0.3481	113.148		
+	0.3482	113.304		
+	0.3483	113.397		
+	0.3484	113.559		
+	0.3485	113.658		
+	0.3486	113.571		
+	0.3487	113.484		
+	0.3488	113.105		
+	0.3489	112.377		
+	0.349	111.22		
+	0.3491	109.715		
+	0.3492	107.569		
+	0.3493	104.403		
+	0.3494	100.235		
+	0.3495	94.369		
+	0.3496	85.257		
+	0.3497	76.94		
+	0.3498	70.291		
+	0.3499	64.021		
+	0.35	58.18		
+	0.3501	53.017		
+	0.3502	48.016		
+	0.3503	43.27		
+	0.3504	38.841		
+	0.3505	34.854		
+	0.3506	30.798		
+	0.3507	27.141		
+	0.3508	23.701		
+	0.3509	20.392		
+	0.351	17.226		
+	0.3511	14.476		
+	0.3512	11.92		
+	0.3513	9.369		
+	0.3514	7.236		
+	0.3515	5.444		
+	0.3516	3.659		
+	0.3517	2.179		
+	0.3518	1.115		
+	0.3519	0.132		
+	0.352	-0.764		
+	0.3521	-1.28		
+	0.3522	-1.777		
+	0.3523	-2.194		
+	0.3524	-2.431		
+	0.3525	-2.487		
+	0.3526	-2.729		
+	0.3527	-2.791		
+	0.3528	-2.717		
+	0.3529	-2.71		
+	0.353	-2.785		
+	0.3531	-2.661		
+	0.3532	-2.599		
+	0.3533	-2.623		
+	0.3534	-2.574		
+	0.3535	-2.424		
+	0.3536	-2.35		
+	0.3537	-2.256		
+	0.3538	-2.151		
+	0.3539	-2.138		
+	0.354	-2.12		
+	0.3541	-2.026		
+	0.3542	-1.945		
+	0.3543	-1.921		
+	0.3544	-1.889		
+	0.3545	-1.809		
+	0.3546	-1.939		
+	0.3547	-1.933		
+	0.3548	-1.771		
+	0.3549	-1.74		
+	0.355	-1.858		
+	0.3551	-1.697		
+	0.3552	-1.591		
+	0.3553	-1.56		
+	0.3554	-1.522		
+	0.3555	-1.274		
+	0.3556	-1.386		
+	0.3557	-1.305		
+	0.3558	-1.243		
+	0.3559	-1.149		
+	0.356	-1.174		
+	0.3561	-0.95		
+	0.3562	-0.963		
+	0.3563	-0.95		
+	0.3564	-0.863		
+	0.3565	-0.689		
+	0.3566	-0.645		
+	0.3567	-0.652		
+	0.3568	-0.502		
+	0.3569	-0.39		
+	0.357	-0.359		
+	0.3571	-0.247		
+	0.3572	-0.117		
+	0.3573	-0.104		
+	0.3574	-0.03		
+	0.3575	0.014		
+	0.3576	0.039		
+	0.3577	-0.054		
+	0.3578	0.026		
+	0.3579	-0.005		
+	0.358	-0.086		
+	0.3581	0.132		
+	0.3582	0.257		
+	0.3583	0.592		
+	0.3584	1.152		
+	0.3585	2.098		
+	0.3586	3.367		
+	0.3587	5.283		
+	0.3588	8.075		
+	0.3589	10.937		
+	0.359	14.19		
+	0.3591	17.891		
+	0.3592	21.99		
+	0.3593	26.164		
+	0.3594	30.755		
+	0.3595	35.675		
+	0.3596	40.769		
+	0.3597	46.243		
+	0.3598	51.904		
+	0.3599	57.763		
+	0.36	63.591		
+	0.3601	69.513		
+	0.3602	75.478		
+	0.3603	81.046		
+	0.3604	86.159		
+	0.3605	90.706		
+	0.3606	93.922		
+	0.3607	96.447		
+	0.3608	98.357		
+	0.3609	99.843		
+	0.361	100.727		
+	0.3611	101.448		
+	0.3612	102.145		
+	0.3613	102.524		
+	0.3614	103.04		
+	0.3615	103.718		
+	0.3616	104.266		
+	0.3617	104.875		
+	0.3618	105.84		
+	0.3619	106.717		
+	0.362	107.432		
+	0.3621	108.154		
+	0.3622	108.863		
+	0.3623	109.429		
+	0.3624	109.933		
+	0.3625	110.455		
+	0.3626	110.872		
+	0.3627	111.04		
+	0.3628	111.313		
+	0.3629	111.568		
+	0.363	111.68		
+	0.3631	111.799		
+	0.3632	111.96		
+	0.3633	111.998		
+	0.3634	112.035		
+	0.3635	112.153		
+	0.3636	112.246		
+	0.3637	112.321		
+	0.3638	112.483		
+	0.3639	112.502		
+	0.364	112.551		
+	0.3641	112.638		
+	0.3642	112.893		
+	0.3643	112.962		
+	0.3644	113.024		
+	0.3645	113.248		
+	0.3646	113.441		
+	0.3647	113.522		
+	0.3648	113.658		
+	0.3649	113.683		
+	0.365	113.503		
+	0.3651	113.242		
+	0.3652	112.912		
+	0.3653	112.166		
+	0.3654	110.872		
+	0.3655	109.248		
+	0.3656	106.773		
+	0.3657	103.463		
+	0.3658	98.966		
+	0.3659	92.242		
+	0.366	83.036		
+	0.3661	75.161		
+	0.3662	68.729		
+	0.3663	62.69		
+	0.3664	56.992		
+	0.3665	51.754		
+	0.3666	46.896		
+	0.3667	42.138		
+	0.3668	37.808		
+	0.3669	33.883		
+	0.367	29.977		
+	0.3671	26.382		
+	0.3672	22.936		
+	0.3673	19.776		
+	0.3674	16.728		
+	0.3675	13.991		
+	0.3676	11.459		
+	0.3677	9.033		
+	0.3678	6.9		
+	0.3679	5.065		
+	0.368	3.416		
+	0.3681	1.998		
+	0.3682	0.816		
+	0.3683	-0.092		
+	0.3684	-0.931		
+	0.3685	-1.479		
+	0.3686	-1.871		
+	0.3687	-2.269		
+	0.3688	-2.468		
+	0.3689	-2.549		
+	0.369	-2.648		
+	0.3691	-2.692		
+	0.3692	-2.592		
+	0.3693	-2.667		
+	0.3694	-2.667		
+	0.3695	-2.692		
+	0.3696	-2.567		
+	0.3697	-2.468		
+	0.3698	-2.505		
+	0.3699	-2.462		
+	0.37	-2.418		
+	0.3701	-2.381		
+	0.3702	-2.244		
+	0.3703	-2.12		
+	0.3704	-2.07		
+	0.3705	-2.039		
+	0.3706	-1.939		
+	0.3707	-1.877		
+	0.3708	-1.939		
+	0.3709	-1.777		
+	0.371	-1.815		
+	0.3711	-1.802		
+	0.3712	-1.79		
+	0.3713	-1.777		
+	0.3714	-1.703		
+	0.3715	-1.728		
+	0.3716	-1.641		
+	0.3717	-1.634		
+	0.3718	-1.628		
+	0.3719	-1.392		
+	0.372	-1.305		
+	0.3721	-1.249		
+	0.3722	-1.28		
+	0.3723	-1.05		
+	0.3724	-0.987		
+	0.3725	-0.907		
+	0.3726	-0.851		
+	0.3727	-0.826		
+	0.3728	-0.832		
+	0.3729	-0.683		
+	0.373	-0.633		
+	0.3731	-0.533		
+	0.3732	-0.459		
+	0.3733	-0.378		
+	0.3734	-0.309		
+	0.3735	-0.291		
+	0.3736	-0.092		
+	0.3737	-0.117		
+	0.3738	-0.042		
+	0.3739	0.026		
+	0.374	0.07		
+	0.3741	0.051		
+	0.3742	0.138		
+	0.3743	0.12		
+	0.3744	0.145		
+	0.3745	0.163		
+	0.3746	0.437		
+	0.3747	0.866		
+	0.3748	1.414		
+	0.3749	2.371		
+	0.375	3.908		
+	0.3751	6.085		
+	0.3752	8.853		
+	0.3753	11.969		
+	0.3754	15.316		
+	0.3755	19.166		
+	0.3756	23.253		
+	0.3757	27.607		
+	0.3758	32.235		
+	0.3759	37.255		
+	0.376	42.474		
+	0.3761	47.96		
+	0.3762	53.651		
+	0.3763	59.48		
+	0.3764	65.358		
+	0.3765	71.093		
+	0.3766	76.89		
+	0.3767	82.439		
+	0.3768	87.365		
+	0.3769	91.527		
+	0.377	94.668		
+	0.3771	96.988		
+	0.3772	98.674		
+	0.3773	100.061		
+	0.3774	100.95		
+	0.3775	101.604		
+	0.3776	102.232		
+	0.3777	102.773		
+	0.3778	103.24		
+	0.3779	103.762		
+	0.378	104.465		
+	0.3781	105.168		
+	0.3782	105.871		
+	0.3783	106.779		
+	0.3784	107.5		
+	0.3785	108.203		
+	0.3786	108.863		
+	0.3787	109.534		
+	0.3788	110.038		
+	0.3789	110.443		
+	0.379	110.785		
+	0.3791	111.108		
+	0.3792	111.425		
+	0.3793	111.618		
+	0.3794	111.799		
+	0.3795	111.861		
+	0.3796	111.917		
+	0.3797	112.097		
+	0.3798	112.035		
+	0.3799	112.041		
+	0.38	112.172		
+	0.3801	112.24		
+	0.3802	112.315		
+	0.3803	112.446		
+	0.3804	112.595		
+	0.3805	112.669		
+	0.3806	112.806		
+	0.3807	112.999		
+	0.3808	113.155		
+	0.3809	113.291		
+	0.381	113.59		
+	0.3811	113.652		
+	0.3812	113.584		
+	0.3813	113.683		
+	0.3814	113.615		
+	0.3815	113.192		
+	0.3816	112.669		
+	0.3817	111.805		
+	0.3818	110.461		
+	0.3819	108.57		
+	0.382	106.132		
+	0.3821	102.63		
+	0.3822	97.66		
+	0.3823	90.227		
+	0.3824	81.307		
+	0.3825	73.886		
+	0.3826	67.467		
+	0.3827	61.576		
+	0.3828	55.978		
+	0.3829	50.803		
+	0.383	45.976		
+	0.3831	41.422		
+	0.3832	37.062		
+	0.3833	33.093		
+	0.3834	29.305		
+	0.3835	25.704		
+	0.3836	22.382		
+	0.3837	19.26		
+	0.3838	16.212		
+	0.3839	13.5		
+	0.384	11.036		
+	0.3841	8.753		
+	0.3842	6.744		
+	0.3843	4.853		
+	0.3844	3.329		
+	0.3845	1.855		
+	0.3846	0.661		
+	0.3847	-0.142		
+	0.3848	-1.019		
+	0.3849	-1.609		
+	0.385	-1.976		
+	0.3851	-2.275		
+	0.3852	-2.561		
+	0.3853	-2.592		
+	0.3854	-2.636		
+	0.3855	-2.661		
+	0.3856	-2.679		
+	0.3857	-2.555		
+	0.3858	-2.543		
+	0.3859	-2.58		
+	0.386	-2.468		
+	0.3861	-2.462		
+	0.3862	-2.53		
+	0.3863	-2.431		
+	0.3864	-2.281		
+	0.3865	-2.343		
+	0.3866	-2.288		
+	0.3867	-2.207		
+	0.3868	-2.144		
+	0.3869	-2.07		
+	0.387	-1.964		
+	0.3871	-1.827		
+	0.3872	-1.908		
+	0.3873	-1.802		
+	0.3874	-1.634		
+	0.3875	-1.684		
+	0.3876	-1.728		
+	0.3877	-1.634		
+	0.3878	-1.684		
+	0.3879	-1.703		
+	0.388	-1.609		
+	0.3881	-1.485		
+	0.3882	-1.541		
+	0.3883	-1.485		
+	0.3884	-1.354		
+	0.3885	-1.342		
+	0.3886	-1.267		
+	0.3887	-1.019		
+	0.3888	-0.95		
+	0.3889	-0.981		
+	0.389	-0.857		
+	0.3891	-0.658		
+	0.3892	-0.633		
+	0.3893	-0.614		
+	0.3894	-0.477		
+	0.3895	-0.49		
+	0.3896	-0.502		
+	0.3897	-0.285		
+	0.3898	-0.229		
+	0.3899	-0.297		
+	0.39	-0.117		
+	0.3901	-0.061		
+	0.3902	-0.079		
+	0.3903	0.014		
+	0.3904	0.176		
+	0.3905	0.107		
+	0.3906	0.002		
+	0.3907	0.244		
+	0.3908	0.275		
+	0.3909	0.294		
+	0.391	0.586		
+	0.3911	1.078		
+	0.3912	1.582		
+	0.3913	2.608		
+	0.3914	4.231		
+	0.3915	6.489		
+	0.3916	9.145		
+	0.3917	12.311		
+	0.3918	15.751		
+	0.3919	19.533		
+	0.392	23.726		
+	0.3921	28.204		
+	0.3922	32.789		
+	0.3923	37.821		
+	0.3924	43.22		
+	0.3925	48.719		
+	0.3926	54.261		
+	0.3927	60.158		
+	0.3928	65.968		
+	0.3929	71.709		
+	0.393	77.432		
+	0.3931	83.024		
+	0.3932	87.745		
+	0.3933	91.614		
+	0.3934	94.73		
+	0.3935	96.963		
+	0.3936	98.637		
+	0.3937	100.024		
+	0.3938	100.957		
+	0.3939	101.529		
+	0.394	102.139		
+	0.3941	102.736		
+	0.3942	103.296		
+	0.3943	103.756		
+	0.3944	104.564		
+	0.3945	105.168		
+	0.3946	105.858		
+	0.3947	106.773		
+	0.3948	107.55		
+	0.3949	108.079		
+	0.395	108.763		
+	0.3951	109.354		
+	0.3952	109.845		
+	0.3953	110.206		
+	0.3954	110.704		
+	0.3955	111.034		
+	0.3956	111.208		
+	0.3957	111.568		
+	0.3958	111.805		
+	0.3959	111.855		
+	0.396	111.979		
+	0.3961	112.06		
+	0.3962	112.004		
+	0.3963	112.016		
+	0.3964	112.209		
+	0.3965	112.166		
+	0.3966	112.135		
+	0.3967	112.253		
+	0.3968	112.458		
+	0.3969	112.446		
+	0.397	112.657		
+	0.3971	112.949		
+	0.3972	113.03		
+	0.3973	113.211		
+	0.3974	113.478		
+	0.3975	113.646		
+	0.3976	113.615		
+	0.3977	113.652		
+	0.3978	113.503		
+	0.3979	113.148		
+	0.398	112.427		
+	0.3981	111.73		
+	0.3982	110.188		
+	0.3983	108.253		
+	0.3984	105.703		
+	0.3985	102.257		
+	0.3986	97.262		
+	0.3987	89.654		
+	0.3988	80.934		
+	0.3989	73.42		
+	0.399	67.143		
+	0.3991	61.445		
+	0.3992	55.853		
+	0.3993	50.647		
+	0.3994	45.864		
+	0.3995	41.248		
+	0.3996	36.844		
+	0.3997	32.975		
+	0.3998	29.231		
+	0.3999	25.449		
+	0.4	22.121		
+	0.4001	19.129		
+	0.4002	16.143		
+	0.4003	13.369		
+	0.4004	10.949		
+	0.4005	8.797		
+	0.4006	6.614		
+	0.4007	4.835		
+	0.4008	3.348		
+	0.4009	1.899		
+	0.401	0.785		
+	0.4011	-0.148		
+	0.4012	-0.944		
+	0.4013	-1.597		
+	0.4014	-1.927		
+	0.4015	-2.244		
+	0.4016	-2.679		
+	0.4017	-2.686		
+	0.4018	-2.661		
+	0.4019	-2.717		
+	0.402	-2.723		
+	0.4021	-2.549		
+	0.4022	-2.561		
+	0.4023	-2.605		
+	0.4024	-2.462		
+	0.4025	-2.337		
+	0.4026	-2.424		
+	0.4027	-2.325		
+	0.4028	-2.194		
+	0.4029	-2.238		
+	0.403	-2.281		
+	0.4031	-2.095		
+	0.4032	-2.151		
+	0.4033	-2.169		
+	0.4034	-1.995		
+	0.4035	-1.889		
+	0.4036	-1.896		
+	0.4037	-1.858		
+	0.4038	-1.616		
+	0.4039	-1.672		
+	0.404	-1.659		
+	0.4041	-1.498		
+	0.4042	-1.466		
+	0.4043	-1.609		
+	0.4044	-1.491		
+	0.4045	-1.41		
+	0.4046	-1.516		
+	0.4047	-1.485		
+	0.4048	-1.261		
+	0.4049	-1.354		
+	0.405	-1.305		
+	0.4051	-1.093		
+	0.4052	-0.95		
+	0.4053	-0.907		
+	0.4054	-0.77		
+	0.4055	-0.558		
+	0.4056	-0.583		
+	0.4057	-0.564		
+	0.4058	-0.359		
+	0.4059	-0.316		
+	0.406	-0.39		
+	0.4061	-0.272		
+	0.4062	-0.185		
+	0.4063	-0.26		
+	0.4064	-0.098		
+	0.4065	0.014		
+	0.4066	-0.086		
+	0.4067	-0.086		
+	0.4068	0.114		
+	0.4069	0.107		
+	0.407	0.002		
+	0.4071	0.294		
+	0.4072	0.294		
+	0.4073	0.319		
+	0.4074	0.692		
+	0.4075	1.264		
+	0.4076	1.855		
+	0.4077	2.906		
+	0.4078	4.692		
+	0.4079	7.074		
+	0.408	9.693		
+	0.4081	12.996		
+	0.4082	16.454		
+	0.4083	20.224		
+	0.4084	24.447		
+	0.4085	28.951		
+	0.4086	33.566		
+	0.4087	38.611		
+	0.4088	44.122		
+	0.4089	49.583		
+	0.409	55.194		
+	0.4091	61.066		
+	0.4092	66.963		
+	0.4093	72.574		
+	0.4094	78.284		
+	0.4095	83.615		
+	0.4096	88.218		
+	0.4097	91.9		
+	0.4098	94.898		
+	0.4099	96.976		
+	0.41	98.5		
+	0.4101	99.793		
+	0.4102	100.739		
+	0.4103	101.305		
+	0.4104	101.971		
+	0.4105	102.605		
+	0.4106	103.022		
+	0.4107	103.712		
+	0.4108	104.484		
+	0.4109	105.205		
+	0.411	105.877		
+	0.4111	106.704		
+	0.4112	107.401		
+	0.4113	107.948		
+	0.4114	108.601		
+	0.4115	109.286		
+	0.4116	109.653		
+	0.4117	109.933		
+	0.4118	110.436		
+	0.4119	110.754		
+	0.412	110.996		
+	0.4121	111.351		
+	0.4122	111.581		
+	0.4123	111.6		
+	0.4124	111.761		
+	0.4125	111.929		
+	0.4126	111.867		
+	0.4127	111.848		
+	0.4128	111.935		
+	0.4129	112.004		
+	0.413	111.917		
+	0.4131	112.066		
+	0.4132	112.178		
+	0.4133	112.215		
+	0.4134	112.296		
+	0.4135	112.607		
+	0.4136	112.806		
+	0.4137	112.937		
+	0.4138	113.279		
+	0.4139	113.366		
+	0.414	113.291		
+	0.4141	113.397		
+	0.4142	113.229		
+	0.4143	112.781		
+	0.4144	112.122		
+	0.4145	111.201		
+	0.4146	109.696		
+	0.4147	107.606		
+	0.4148	104.907		
+	0.4149	101.162		
+	0.415	95.9		
+	0.4151	87.813		
+	0.4152	79.291		
+	0.4153	72.132		
+	0.4154	66.017		
+	0.4155	60.326		
+	0.4156	54.889		
+	0.4157	49.776		
+	0.4158	44.993		
+	0.4159	40.452		
+	0.416	36.197		
+	0.4161	32.279		
+	0.4162	28.584		
+	0.4163	24.97		
+	0.4164	21.567		
+	0.4165	18.538		
+	0.4166	15.633		
+	0.4167	12.772		
+	0.4168	10.483		
+	0.4169	8.349		
+	0.417	6.259		
+	0.4171	4.586		
+	0.4172	3.056		
+	0.4173	1.725		
+	0.4174	0.636		
+	0.4175	-0.229		
+	0.4176	-0.95		
+	0.4177	-1.634		
+	0.4178	-2.07		
+	0.4179	-2.312		
+	0.418	-2.605		
+	0.4181	-2.698		
+	0.4182	-2.71		
+	0.4183	-2.76		
+	0.4184	-2.829		
+	0.4185	-2.636		
+	0.4186	-2.617		
+	0.4187	-2.549		
+	0.4188	-2.381		
+	0.4189	-2.368		
+	0.419	-2.387		
+	0.4191	-2.312		
+	0.4192	-2.213		
+	0.4193	-2.176		
+	0.4194	-2.219		
+	0.4195	-2.132		
+	0.4196	-2.088		
+	0.4197	-2.132		
+	0.4198	-2.02		
+	0.4199	-1.933		
+	0.42	-1.939		
+	0.4201	-1.889		
+	0.4202	-1.734		
+	0.4203	-1.728		
+	0.4204	-1.684		
+	0.4205	-1.535		
+	0.4206	-1.522		
+	0.4207	-1.491		
+	0.4208	-1.41		
+	0.4209	-1.379		
+	0.421	-1.435		
+	0.4211	-1.41		
+	0.4212	-1.323		
+	0.4213	-1.354		
+	0.4214	-1.236		
+	0.4215	-1.124		
+	0.4216	-0.987		
+	0.4217	-1.006		
+	0.4218	-0.888		
+	0.4219	-0.708		
+	0.422	-0.664		
+	0.4221	-0.54		
+	0.4222	-0.428		
+	0.4223	-0.347		
+	0.4224	-0.341		
+	0.4225	-0.197		
+	0.4226	-0.061		
+	0.4227	-0.098		
+	0.4228	-0.11		
+	0.4229	0.008		
+	0.423	-0.005		
+	0.4231	-0.023		
+	0.4232	0.045		
+	0.4233	0.089		
+	0.4234	-0.048		
+	0.4235	0.138		
+	0.4236	0.194		
+	0.4237	0.362		
+	0.4238	0.686		
+	0.4239	1.183		
+	0.424	1.917		
+	0.4241	3.006		
+	0.4242	4.853		
+	0.4243	7.205		
+	0.4244	9.91		
+	0.4245	13.014		
+	0.4246	16.597		
+	0.4247	20.448		
+	0.4248	24.547		
+	0.4249	29.038		
+	0.425	33.722		
+	0.4251	38.679		
+	0.4252	44.141		
+	0.4253	49.614		
+	0.4254	55.331		
+	0.4255	61.134		
+	0.4256	66.919		
+	0.4257	72.654		
+	0.4258	78.284		
+	0.4259	83.639		
+	0.426	88.224		
+	0.4261	91.819		
+	0.4262	94.649		
+	0.4263	96.808		
+	0.4264	98.413		
+	0.4265	99.563		
+	0.4266	100.459		
+	0.4267	101.125		
+	0.4268	101.647		
+	0.4269	102.275		
+	0.427	102.81		
+	0.4271	103.501		
+	0.4272	104.191		
+	0.4273	104.987		
+	0.4274	105.74		
+	0.4275	106.499		
+	0.4276	107.295		
+	0.4277	107.892		
+	0.4278	108.415		
+	0.4279	109.018		
+	0.428	109.472		
+	0.4281	109.833		
+	0.4282	110.138		
+	0.4283	110.486		
+	0.4284	110.735		
+	0.4285	110.978		
+	0.4286	111.251		
+	0.4287	111.425		
+	0.4288	111.6		
+	0.4289	111.674		
+	0.429	111.73		
+	0.4291	111.68		
+	0.4292	111.811		
+	0.4293	111.83		
+	0.4294	111.811		
+	0.4295	111.861		
+	0.4296	111.973		
+	0.4297	112.116		
+	0.4298	112.147		
+	0.4299	112.352		
+	0.43	112.564		
+	0.4301	112.669		
+	0.4302	112.974		
+	0.4303	113.117		
+	0.4304	113.148		
+	0.4305	113.167		
+	0.4306	113.049		
+	0.4307	112.638		
+	0.4308	111.935		
+	0.4309	111.046		
+	0.431	109.584		
+	0.4311	107.413		
+	0.4312	104.714		
+	0.4313	100.988		
+	0.4314	95.763		
+	0.4315	87.633		
+	0.4316	79.018		
+	0.4317	72.014		
+	0.4318	65.762		
+	0.4319	60.065		
+	0.432	54.703		
+	0.4321	49.72		
+	0.4322	44.868		
+	0.4323	40.458		
+	0.4324	36.21		
+	0.4325	32.291		
+	0.4326	28.596		
+	0.4327	25.032		
+	0.4328	21.648		
+	0.4329	18.47		
+	0.433	15.633		
+	0.4331	12.846		
+	0.4332	10.402		
+	0.4333	8.256		
+	0.4334	6.216		
+	0.4335	4.499		
+	0.4336	3.012		
+	0.4337	1.774		
+	0.4338	0.617		
+	0.4339	-0.247		
+	0.434	-0.925		
+	0.4341	-1.535		
+	0.4342	-2.001		
+	0.4343	-2.238		
+	0.4344	-2.48		
+	0.4345	-2.617		
+	0.4346	-2.704		
+	0.4347	-2.673		
+	0.4348	-2.735		
+	0.4349	-2.729		
+	0.435	-2.642		
+	0.4351	-2.648		
+	0.4352	-2.58		
+	0.4353	-2.387		
+	0.4354	-2.406		
+	0.4355	-2.294		
+	0.4356	-2.219		
+	0.4357	-2.151		
+	0.4358	-2.088		
+	0.4359	-2.057		
+	0.436	-2.02		
+	0.4361	-2.045		
+	0.4362	-2.057		
+	0.4363	-1.958		
+	0.4364	-1.871		
+	0.4365	-1.871		
+	0.4366	-1.833		
+	0.4367	-1.765		
+	0.4368	-1.721		
+	0.4369	-1.697		
+	0.437	-1.572		
+	0.4371	-1.473		
+	0.4372	-1.491		
+	0.4373	-1.348		
+	0.4374	-1.373		
+	0.4375	-1.336		
+	0.4376	-1.274		
+	0.4377	-1.174		
+	0.4378	-1.18		
+	0.4379	-1.124		
+	0.438	-1.006		
+	0.4381	-0.931		
+	0.4382	-0.931		
+	0.4383	-0.764		
+	0.4384	-0.714		
+	0.4385	-0.664		
+	0.4386	-0.453		
+	0.4387	-0.322		
+	0.4388	-0.229		
+	0.4389	-0.191		
+	0.439	-0.086		
+	0.4391	0.045		
+	0.4392	-0.042		
+	0.4393	0.082		
+	0.4394	0.051		
+	0.4395	-0.005		
+	0.4396	0.002		
+	0.4397	0.114		
+	0.4398	0.008		
+	0.4399	0.008		
+	0.44	0.163		
+	0.4401	0.331		
+	0.4402	0.648		
+	0.4403	1.227		
+	0.4404	2.104		
+	0.4405	3.23		
+	0.4406	5.127		
+	0.4407	7.628		
+	0.4408	10.433		
+	0.4409	13.668		
+	0.441	17.201		
+	0.4411	21.076		
+	0.4412	25.088		
+	0.4413	29.56		
+	0.4414	34.437		
+	0.4415	39.376		
+	0.4416	44.638		
+	0.4417	50.23		
+	0.4418	55.897		
+	0.4419	61.545		
+	0.442	67.442		
+	0.4421	73.214		
+	0.4422	78.676		
+	0.4423	83.975		
+	0.4424	88.504		
+	0.4425	92.043		
+	0.4426	94.78		
+	0.4427	96.907		
+	0.4428	98.406		
+	0.4429	99.538		
+	0.443	100.378		
+	0.4431	101.137		
+	0.4432	101.548		
+	0.4433	102.157		
+	0.4434	102.748		
+	0.4435	103.364		
+	0.4436	104.048		
+	0.4437	104.931		
+	0.4438	105.709		
+	0.4439	106.399		
+	0.444	107.227		
+	0.4441	107.923		
+	0.4442	108.421		
+	0.4443	108.993		
+	0.4444	109.466		
+	0.4445	109.733		
+	0.4446	109.989		
+	0.4447	110.43		
+	0.4448	110.673		
+	0.4449	110.797		
+	0.445	111.065		
+	0.4451	111.245		
+	0.4452	111.394		
+	0.4453	111.481		
+	0.4454	111.668		
+	0.4455	111.6		
+	0.4456	111.568		
+	0.4457	111.755		
+	0.4458	111.792		
+	0.4459	111.799		
+	0.446	111.973		
+	0.4461	112.091		
+	0.4462	112.023		
+	0.4463	112.203		
+	0.4464	112.489		
+	0.4465	112.576		
+	0.4466	112.707		
+	0.4467	112.962		
+	0.4468	112.931		
+	0.4469	112.875		
+	0.447	112.781		
+	0.4471	112.446		
+	0.4472	111.705		
+	0.4473	110.704		
+	0.4474	109.217		
+	0.4475	107.077		
+	0.4476	104.185		
+	0.4477	100.403		
+	0.4478	94.911		
+	0.4479	86.364		
+	0.448	78.029		
+	0.4481	71.255		
+	0.4482	64.979		
+	0.4483	59.281		
+	0.4484	54.087		
+	0.4485	49.055		
+	0.4486	44.277		
+	0.4487	40.004		
+	0.4488	35.874		
+	0.4489	31.806		
+	0.449	28.155		
+	0.4491	24.74		
+	0.4492	21.368		
+	0.4493	18.19		
+	0.4494	15.484		
+	0.4495	12.678		
+	0.4496	10.11		
+	0.4497	8.051		
+	0.4498	6.06		
+	0.4499	4.275		
+	0.45	2.788		
+	0.4501	1.55		
+	0.4502	0.449		
+	0.4503	-0.453		
+	0.4504	-0.938		
+	0.4505	-1.541		
+	0.4506	-2.039		
+	0.4507	-2.263		
+	0.4508	-2.437		
+	0.4509	-2.636		
+	0.451	-2.648		
+	0.4511	-2.692		
+	0.4512	-2.71		
+	0.4513	-2.798		
+	0.4514	-2.605		
+	0.4515	-2.599		
+	0.4516	-2.623		
+	0.4517	-2.518		
+	0.4518	-2.412		
+	0.4519	-2.387		
+	0.452	-2.238		
+	0.4521	-2.132		
+	0.4522	-2.157		
+	0.4523	-2.132		
+	0.4524	-2.001		
+	0.4525	-1.889		
+	0.4526	-1.983		
+	0.4527	-1.877		
+	0.4528	-1.827		
+	0.4529	-1.908		
+	0.453	-1.833		
+	0.4531	-1.74		
+	0.4532	-1.79		
+	0.4533	-1.815		
+	0.4534	-1.684		
+	0.4535	-1.529		
+	0.4536	-1.616		
+	0.4537	-1.386		
+	0.4538	-1.286		
+	0.4539	-1.429		
+	0.454	-1.286		
+	0.4541	-1.099		
+	0.4542	-1.081		
+	0.4543	-0.994		
+	0.4544	-0.963		
+	0.4545	-0.894		
+	0.4546	-0.931		
+	0.4547	-0.795		
+	0.4548	-0.652		
+	0.4549	-0.658		
+	0.455	-0.614		
+	0.4551	-0.384		
+	0.4552	-0.316		
+	0.4553	-0.297		
+	0.4554	-0.017		
+	0.4555	0.064		
+	0.4556	-0.036		
+	0.4557	0.12		
+	0.4558	0.201		
+	0.4559	0.051		
+	0.456	0.089		
+	0.4561	0.145		
+	0.4562	0.17		
+	0.4563	0.014		
+	0.4564	0.188		
+	0.4565	0.431		
+	0.4566	0.58		
+	0.4567	1.14		
+	0.4568	1.98		
+	0.4569	3.112		
+	0.457	4.878		
+	0.4571	7.509		
+	0.4572	10.178		
+	0.4573	13.245		
+	0.4574	16.89		
+	0.4575	20.715		
+	0.4576	24.802		
+	0.4577	29.2		
+	0.4578	33.946		
+	0.4579	38.86		
+	0.458	44.047		
+	0.4581	49.664		
+	0.4582	55.163		
+	0.4583	60.836		
+	0.4584	66.733		
+	0.4585	72.381		
+	0.4586	77.917		
+	0.4587	83.254		
+	0.4588	87.975		
+	0.4589	91.508		
+	0.459	94.326		
+	0.4591	96.59		
+	0.4592	98.151		
+	0.4593	99.252		
+	0.4594	100.248		
+	0.4595	100.95		
+	0.4596	101.386		
+	0.4597	101.971		
+	0.4598	102.605		
+	0.4599	103.103		
+	0.46	103.768		
+	0.4601	104.62		
+	0.4602	105.441		
+	0.4603	106.107		
+	0.4604	107.009		
+	0.4605	107.724		
+	0.4606	108.234		
+	0.4607	108.8		
+	0.4608	109.36		
+	0.4609	109.715		
+	0.461	109.989		
+	0.4611	110.318		
+	0.4612	110.573		
+	0.4613	110.66		
+	0.4614	110.99		
+	0.4615	111.201		
+	0.4616	111.226		
+	0.4617	111.307		
+	0.4618	111.5		
+	0.4619	111.544		
+	0.462	111.544		
+	0.4621	111.674		
+	0.4622	111.743		
+	0.4623	111.761		
+	0.4624	111.886		
+	0.4625	112.06		
+	0.4626	112.128		
+	0.4627	112.178		
+	0.4628	112.47		
+	0.4629	112.545		
+	0.463	112.57		
+	0.4631	112.9		
+	0.4632	112.887		
+	0.4633	112.819		
+	0.4634	112.663		
+	0.4635	112.458		
+	0.4636	111.73		
+	0.4637	110.772		
+	0.4638	109.441		
+	0.4639	107.395		
+	0.464	104.596		
+	0.4641	101.131		
+	0.4642	95.999		
+	0.4643	87.981		
+	0.4644	79.391		
+	0.4645	72.35		
+	0.4646	66.036		
+	0.4647	60.32		
+	0.4648	54.964		
+	0.4649	49.894		
+	0.465	45.092		
+	0.4651	40.645		
+	0.4652	36.533		
+	0.4653	32.459		
+	0.4654	28.851		
+	0.4655	25.436		
+	0.4656	22.04		
+	0.4657	18.868		
+	0.4658	16.031		
+	0.4659	13.288		
+	0.466	10.744		
+	0.4661	8.579		
+	0.4662	6.508		
+	0.4663	4.623		
+	0.4664	3.124		
+	0.4665	1.874		
+	0.4666	0.611		
+	0.4667	-0.316		
+	0.4668	-0.894		
+	0.4669	-1.498		
+	0.467	-2.026		
+	0.4671	-2.207		
+	0.4672	-2.387		
+	0.4673	-2.549		
+	0.4674	-2.599		
+	0.4675	-2.518		
+	0.4676	-2.648		
+	0.4677	-2.655		
+	0.4678	-2.518		
+	0.4679	-2.536		
+	0.468	-2.63		
+	0.4681	-2.48		
+	0.4682	-2.399		
+	0.4683	-2.449		
+	0.4684	-2.443		
+	0.4685	-2.151		
+	0.4686	-2.219		
+	0.4687	-2.12		
+	0.4688	-1.952		
+	0.4689	-1.983		
+	0.469	-1.958		
+	0.4691	-1.846		
+	0.4692	-1.746		
+	0.4693	-1.79		
+	0.4694	-1.796		
+	0.4695	-1.715		
+	0.4696	-1.784		
+	0.4697	-1.715		
+	0.4698	-1.672		
+	0.4699	-1.628		
+	0.47	-1.603		
+	0.4701	-1.504		
+	0.4702	-1.361		
+	0.4703	-1.404		
+	0.4704	-1.224		
+	0.4705	-1.087		
+	0.4706	-1.093		
+	0.4707	-1.019		
+	0.4708	-0.863		
+	0.4709	-0.813		
+	0.471	-0.776		
+	0.4711	-0.708		
+	0.4712	-0.558		
+	0.4713	-0.664		
+	0.4714	-0.527		
+	0.4715	-0.341		
+	0.4716	-0.372		
+	0.4717	-0.291		
+	0.4718	-0.148		
+	0.4719	-0.067		
+	0.472	0.008		
+	0.4721	0.101		
+	0.4722	0.157		
+	0.4723	0.157		
+	0.4724	0.176		
+	0.4725	0.306		
+	0.4726	0.225		
+	0.4727	0.176		
+	0.4728	0.294		
+	0.4729	0.418		
+	0.473	0.53		
+	0.4731	0.207		
+	0.4732	0.81		
+	0.4733	1.805		
+	0.4734	3.267		
+	0.4735	5.32		
+	0.4736	8.026		
+	0.4737	11.385		
+	0.4738	15.129		
+	0.4739	19.123		
+	0.474	23.508		
+	0.4741	28.534		
+	0.4742	33.622		
+	0.4743	39.071		
+	0.4744	45.211		
+	0.4745	51.493		
+	0.4746	57.943		
+	0.4747	64.661		
+	0.4748	71.448		
+	0.4749	77.998		
+	0.475	84.286		
+	0.4751	89.773		
+	0.4752	93.803		
+	0.4753	96.739		
+	0.4754	99.004		
+	0.4755	100.49		
+	0.4756	101.38		
+	0.4757	102.039		
+	0.4758	102.593		
+	0.4759	102.922		
+	0.476	103.482		
+	0.4761	104.135		
+	0.4762	104.745		
+	0.4763	105.473		
+	0.4764	106.381		
+	0.4765	107.245		
+	0.4766	107.874		
+	0.4767	108.72		
+	0.4768	109.366		
+	0.4769	109.796		
+	0.477	110.237		
+	0.4771	110.685		
+	0.4772	111.009		
+	0.4773	111.096		
+	0.4774	111.345		
+	0.4775	111.519		
+	0.4776	111.5		
+	0.4777	111.631		
+	0.4778	111.824		
+	0.4779	111.656		
+	0.478	111.724		
+	0.4781	111.805		
+	0.4782	111.792		
+	0.4783	111.736		
+	0.4784	111.83		
+	0.4785	111.836		
+	0.4786	111.699		
+	0.4787	111.749		
+	0.4788	111.979		
+	0.4789	111.898		
+	0.479	112.004		
+	0.4791	112.315		
+	0.4792	112.352		
+	0.4793	112.396		
+	0.4794	112.526		
+	0.4795	112.483		
+	0.4796	112.29		
+	0.4797	111.867		
+	0.4798	111.369		
+	0.4799	110.256		
+	0.48	108.626		
+	0.4801	106.511		
+	0.4802	103.246		
+	0.4803	98.587		
+	0.4804	91.962		
+	0.4805	82.29		
+	0.4806	73.42		
+	0.4807	66.384		
+	0.4808	60.145		
+	0.4809	54.112		
+	0.481	48.576		
+	0.4811	43.494		
+	0.4812	38.692		
+	0.4813	34.089		
+	0.4814	30.058		
+	0.4815	26.326		
+	0.4816	22.625		
+	0.4817	19.309		
+	0.4818	16.33		
+	0.4819	13.468		
+	0.482	10.738		
+	0.4821	8.498		
+	0.4822	6.365		
+	0.4823	4.399		
+	0.4824	2.782		
+	0.4825	1.407		
+	0.4826	0.194		
+	0.4827	-0.757		
+	0.4828	-1.46		
+	0.4829	-2.064		
+	0.483	-2.599		
+	0.4831	-2.804		
+	0.4832	-2.99		
+	0.4833	-3.158		
+	0.4834	-3.127		
+	0.4835	-2.99		
+	0.4836	-3.127		
+	0.4837	-3.077		
+	0.4838	-2.922		
+	0.4839	-2.941		
+	0.484	-2.947		
+	0.4841	-2.866		
+	0.4842	-2.791		
+	0.4843	-2.866		
+	0.4844	-2.717		
+	0.4845	-2.623		
+	0.4846	-2.655		
+	0.4847	-2.636		
+	0.4848	-2.431		
+	0.4849	-2.381		
+	0.485	-2.381		
+	0.4851	-2.269		
+	0.4852	-2.132		
+	0.4853	-2.138		
+	0.4854	-2.182		
+	0.4855	-2.057		
+	0.4856	-2.076		
+	0.4857	-2.207		
+	0.4858	-2.076		
+	0.4859	-2.032		
+	0.486	-2.032		
+	0.4861	-1.952		
+	0.4862	-1.952		
+	0.4863	-2.02		
+	0.4864	-1.914		
+	0.4865	-1.678		
+	0.4866	-1.703		
+	0.4867	-1.585		
+	0.4868	-1.529		
+	0.4869	-1.442		
+	0.487	-1.442		
+	0.4871	-1.336		
+	0.4872	-1.205		
+	0.4873	-1.274		
+	0.4874	-1.23		
+	0.4875	-1.081		
+	0.4876	-1.131		
+	0.4877	-1.081		
+	0.4878	-1.019		
+	0.4879	-0.931		
+	0.488	-0.963		
+	0.4881	-0.857		
+	0.4882	-0.72		
+	0.4883	-0.72		
+	0.4884	-0.676		
+	0.4885	-0.515		
+	0.4886	-0.521		
+	0.4887	-0.589		
+	0.4888	-0.471		
+	0.4889	-0.477		
+	0.489	-0.496		
+	0.4891	-0.372		
+	0.4892	-0.079		
+	0.4893	0.188		
+	0.4894	0.841		
+	0.4895	1.924		
+	0.4896	3.292		
+	0.4897	5.382		
+	0.4898	8.393		
+	0.4899	11.633		
+	0.49	15.366		
+	0.4901	19.515		
+	0.4902	24.118		
+	0.4903	28.926		
+	0.4904	34.114		
+	0.4905	39.743		
+	0.4906	45.77		
+	0.4907	51.879		
+	0.4908	58.385		
+	0.4909	64.979		
+	0.491	71.616		
+	0.4911	78.122		
+	0.4912	84.429		
+	0.4913	89.605		
+	0.4914	93.722		
+	0.4915	96.721		
+	0.4916	98.929		
+	0.4917	100.403		
+	0.4918	101.367		
+	0.4919	102.058		
+	0.492	102.58		
+	0.4921	103.04		
+	0.4922	103.575		
+	0.4923	104.073		
+	0.4924	104.739		
+	0.4925	105.553		
+	0.4926	106.3		
+	0.4927	107.084		
+	0.4928	107.843		
+	0.4929	108.589		
+	0.493	109.074		
+	0.4931	109.646		
+	0.4932	110.256		
+	0.4933	110.573		
+	0.4934	110.841		
+	0.4935	111.164		
+	0.4936	111.394		
+	0.4937	111.432		
+	0.4938	111.624		
+	0.4939	111.705		
+	0.494	111.712		
+	0.4941	111.705		
+	0.4942	111.805		
+	0.4943	111.755		
+	0.4944	111.755		
+	0.4945	111.792		
+	0.4946	111.712		
+	0.4947	111.587		
+	0.4948	111.593		
+	0.4949	111.792		
+	0.495	111.799		
+	0.4951	111.935		
+	0.4952	112.103		
+	0.4953	112.309		
+	0.4954	112.421		
+	0.4955	112.595		
+	0.4956	112.613		
+	0.4957	112.539		
+	0.4958	112.358		
+	0.4959	111.979		
+	0.496	111.276		
+	0.4961	110.206		
+	0.4962	108.626		
+	0.4963	106.325		
+	0.4964	103.04		
+	0.4965	98.531		
+	0.4966	91.937		
+	0.4967	82.171		
+	0.4968	73.488		
+	0.4969	66.54		
+	0.497	60.201		
+	0.4971	54.199		
+	0.4972	48.744		
+	0.4973	43.618		
+	0.4974	38.766		
+	0.4975	34.325		
+	0.4976	30.12		
+	0.4977	26.338		
+	0.4978	22.643		
+	0.4979	19.353		
+	0.498	16.205		
+	0.4981	13.363		
+	0.4982	10.844		
+	0.4983	8.573		
+	0.4984	6.415		
+	0.4985	4.598		
+	0.4986	3.012		
+	0.4987	1.55		
+	0.4988	0.381		
+	0.4989	-0.533		
+	0.499	-1.342		
+	0.4991	-2.032		
+	0.4992	-2.431		
+	0.4993	-2.779		
+	0.4994	-3.028		
+	0.4995	-3.14		
+	0.4996	-3.196		
+	0.4997	-3.165		
+	0.4998	-3.165		
+	0.4999	-3.046		
+	0.5	-2.941		
+	0.5001	-2.934		
+	0.5002	-2.922		
+	0.5003	-2.785		
+	0.5004	-2.729		
+	0.5005	-2.692		
+	0.5006	-2.58		
+	0.5007	-2.605		
+	0.5008	-2.536		
+	0.5009	-2.518		
+	0.501	-2.418		
+	0.5011	-2.443		
+	0.5012	-2.362		
+	0.5013	-2.35		
+	0.5014	-2.263		
+	0.5015	-2.25		
+	0.5016	-2.126		
+	0.5017	-2.126		
+	0.5018	-2.12		
+	0.5019	-2.064		
+	0.502	-1.995		
+	0.5021	-2.001		
+	0.5022	-1.933		
+	0.5023	-1.833		
+	0.5024	-1.921		
+	0.5025	-1.883		
+	0.5026	-1.765		
+	0.5027	-1.734		
+	0.5028	-1.753		
+	0.5029	-1.653		
+	0.503	-1.554		
+	0.5031	-1.628		
+	0.5032	-1.485		
+	0.5033	-1.323		
+	0.5034	-1.323		
+	0.5035	-1.298		
+	0.5036	-1.143		
+	0.5037	-0.994		
+	0.5038	-1.037		
+	0.5039	-0.9		
+	0.504	-0.876		
+	0.5041	-0.9		
+	0.5042	-0.9		
+	0.5043	-0.77		
+	0.5044	-0.788		
+	0.5045	-0.77		
+	0.5046	-0.714		
+	0.5047	-0.62		
+	0.5048	-0.701		
+	0.5049	-0.546		
+	0.505	-0.49		
+	0.5051	-0.459		
+	0.5052	-0.428		
+	0.5053	-0.272		
+	0.5054	-0.067		
+	0.5055	0.313		
+	0.5056	0.966		
+	0.5057	1.893		
+	0.5058	3.217		
+	0.5059	5.233		
+	0.506	8.163		
+	0.5061	11.31		
+	0.5062	14.974		
+	0.5063	19.085		
+	0.5064	23.496		
+	0.5065	28.248		
+	0.5066	33.535		
+	0.5067	39.04		
+	0.5068	44.937		
+	0.5069	51.12		
+	0.507	57.651		
+	0.5071	64.182		
+	0.5072	70.745		
+	0.5073	77.289		
+	0.5074	83.552		
+	0.5075	88.821		
+	0.5076	93.057		
+	0.5077	96.223		
+	0.5078	98.413		
+	0.5079	99.961		
+	0.508	101.069		
+	0.5081	101.703		
+	0.5082	102.25		
+	0.5083	102.823		
+	0.5084	103.37		
+	0.5085	103.886		
+	0.5086	104.602		
+	0.5087	105.466		
+	0.5088	106.144		
+	0.5089	106.941		
+	0.509	107.737		
+	0.5091	108.353		
+	0.5092	108.937		
+	0.5093	109.578		
+	0.5094	110.094		
+	0.5095	110.331		
+	0.5096	110.648		
+	0.5097	110.953		
+	0.5098	111.096		
+	0.5099	111.351		
+	0.51	111.5		
+	0.5101	111.649		
+	0.5102	111.662		
+	0.5103	111.712		
+	0.5104	111.768		
+	0.5105	111.755		
+	0.5106	111.805		
+	0.5107	111.768		
+	0.5108	111.687		
+	0.5109	111.55		
+	0.511	111.693		
+	0.5111	111.593		
+	0.5112	111.612		
+	0.5113	111.768		
+	0.5114	111.985		
+	0.5115	112.097		
+	0.5116	112.296		
+	0.5117	112.489		
+	0.5118	112.526		
+	0.5119	112.502		
+	0.512	112.402		
+	0.5121	112.147		
+	0.5122	111.376		
+	0.5123	110.455		
+	0.5124	108.987		
+	0.5125	106.623		
+	0.5126	103.607		
+	0.5127	99.377		
+	0.5128	93.113		
+	0.5129	83.615		
+	0.513	74.744		
+	0.5131	67.572		
+	0.5132	61.141		
+	0.5133	55.194		
+	0.5134	49.789		
+	0.5135	44.489		
+	0.5136	39.631		
+	0.5137	35.277		
+	0.5138	31.003		
+	0.5139	27.035		
+	0.514	23.502		
+	0.5141	20.012		
+	0.5142	16.809		
+	0.5143	13.935		
+	0.5144	11.341		
+	0.5145	8.828		
+	0.5146	6.701		
+	0.5147	4.884		
+	0.5148	3.168		
+	0.5149	1.749		
+	0.515	0.611		
+	0.5151	-0.328		
+	0.5152	-1.311		
+	0.5153	-1.765		
+	0.5154	-2.219		
+	0.5155	-2.642		
+	0.5156	-2.872		
+	0.5157	-2.934		
+	0.5158	-3.152		
+	0.5159	-3.239		
+	0.516	-3.096		
+	0.5161	-3.04		
+	0.5162	-3.146		
+	0.5163	-2.997		
+	0.5164	-2.953		
+	0.5165	-2.947		
+	0.5166	-2.866		
+	0.5167	-2.655		
+	0.5168	-2.592		
+	0.5169	-2.648		
+	0.517	-2.368		
+	0.5171	-2.362		
+	0.5172	-2.393		
+	0.5173	-2.343		
+	0.5174	-2.232		
+	0.5175	-2.331		
+	0.5176	-2.3		
+	0.5177	-2.163		
+	0.5178	-2.188		
+	0.5179	-2.294		
+	0.518	-2.2		
+	0.5181	-2.082		
+	0.5182	-2.107		
+	0.5183	-2.001		
+	0.5184	-1.852		
+	0.5185	-1.939		
+	0.5186	-1.883		
+	0.5187	-1.715		
+	0.5188	-1.672		
+	0.5189	-1.784		
+	0.519	-1.585		
+	0.5191	-1.566		
+	0.5192	-1.585		
+	0.5193	-1.572		
+	0.5194	-1.354		
+	0.5195	-1.448		
+	0.5196	-1.473		
+	0.5197	-1.23		
+	0.5198	-1.131		
+	0.5199	-1.187		
+	0.52	-0.963		
+	0.5201	-0.801		
+	0.5202	-0.931		
+	0.5203	-0.838		
+	0.5204	-0.664		
+	0.5205	-0.708		
+	0.5206	-0.745		
+	0.5207	-0.627		
+	0.5208	-0.62		
+	0.5209	-0.708		
+	0.521	-0.571		
+	0.5211	-0.552		
+	0.5212	-0.645		
+	0.5213	-0.67		
+	0.5214	-0.465		
+	0.5215	-0.39		
+	0.5216	-0.21		
+	0.5217	0.356		
+	0.5218	0.991		
+	0.5219	1.861		
+	0.522	3.242		
+	0.5221	5.301		
+	0.5222	8.026		
+	0.5223	11.173		
+	0.5224	14.787		
+	0.5225	18.743		
+	0.5226	23.066		
+	0.5227	27.887		
+	0.5228	33		
+	0.5229	38.343		
+	0.523	44.203		
+	0.5231	50.454		
+	0.5232	56.718		
+	0.5233	63.224		
+	0.5234	69.924		
+	0.5235	76.306		
+	0.5236	82.563		
+	0.5237	88.174		
+	0.5238	92.522		
+	0.5239	95.682		
+	0.524	98.046		
+	0.5241	99.793		
+	0.5242	100.764		
+	0.5243	101.386		
+	0.5244	102.126		
+	0.5245	102.543		
+	0.5246	102.96		
+	0.5247	103.656		
+	0.5248	104.353		
+	0.5249	104.963		
+	0.525	105.889		
+	0.5251	106.841		
+	0.5252	107.476		
+	0.5253	108.185		
+	0.5254	108.869		
+	0.5255	109.435		
+	0.5256	109.827		
+	0.5257	110.268		
+	0.5258	110.648		
+	0.5259	110.754		
+	0.526	111.04		
+	0.5261	111.295		
+	0.5262	111.301		
+	0.5263	111.295		
+	0.5264	111.562		
+	0.5265	111.568		
+	0.5266	111.519		
+	0.5267	111.755		
+	0.5268	111.73		
+	0.5269	111.643		
+	0.527	111.624		
+	0.5271	111.656		
+	0.5272	111.531		
+	0.5273	111.581		
+	0.5274	111.631		
+	0.5275	111.743		
+	0.5276	111.736		
+	0.5277	112.035		
+	0.5278	112.159		
+	0.5279	112.246		
+	0.528	112.246		
+	0.5281	112.377		
+	0.5282	112.222		
+	0.5283	111.898		
+	0.5284	111.425		
+	0.5285	110.536		
+	0.5286	108.968		
+	0.5287	107.028		
+	0.5288	104.135		
+	0.5289	99.974		
+	0.529	94.121		
+	0.5291	85.182		
+	0.5292	75.814		
+	0.5293	68.418		
+	0.5294	62.123		
+	0.5295	56.046		
+	0.5296	50.38		
+	0.5297	45.223		
+	0.5298	40.371		
+	0.5299	35.737		
+	0.53	31.601		
+	0.5301	27.806		
+	0.5302	23.981		
+	0.5303	20.497		
+	0.5304	17.499		
+	0.5305	14.569		
+	0.5306	11.783		
+	0.5307	9.357		
+	0.5308	7.242		
+	0.5309	5.146		
+	0.531	3.441		
+	0.5311	2.06		
+	0.5312	0.754		
+	0.5313	-0.39		
+	0.5314	-1.131		
+	0.5315	-1.765		
+	0.5316	-2.3		
+	0.5317	-2.561		
+	0.5318	-2.692		
+	0.5319	-2.978		
+	0.532	-3.09		
+	0.5321	-2.941		
+	0.5322	-2.978		
+	0.5323	-3.084		
+	0.5324	-2.953		
+	0.5325	-2.966		
+	0.5326	-3.077		
+	0.5327	-2.941		
+	0.5328	-2.822		
+	0.5329	-2.835		
+	0.533	-2.754		
+	0.5331	-2.561		
+	0.5332	-2.474		
+	0.5333	-2.53		
+	0.5334	-2.35		
+	0.5335	-2.269		
+	0.5336	-2.325		
+	0.5337	-2.232		
+	0.5338	-2.057		
+	0.5339	-2.163		
+	0.534	-2.225		
+	0.5341	-2.088		
+	0.5342	-2.157		
+	0.5343	-2.194		
+	0.5344	-2.07		
+	0.5345	-2.001		
+	0.5346	-2.07		
+	0.5347	-2.001		
+	0.5348	-1.871		
+	0.5349	-1.846		
+	0.535	-1.784		
+	0.5351	-1.622		
+	0.5352	-1.597		
+	0.5353	-1.622		
+	0.5354	-1.442		
+	0.5355	-1.33		
+	0.5356	-1.423		
+	0.5357	-1.361		
+	0.5358	-1.211		
+	0.5359	-1.298		
+	0.536	-1.236		
+	0.5361	-1.062		
+	0.5362	-1.106		
+	0.5363	-1.099		
+	0.5364	-0.907		
+	0.5365	-0.869		
+	0.5366	-0.813		
+	0.5367	-0.745		
+	0.5368	-0.589		
+	0.5369	-0.645		
+	0.537	-0.583		
+	0.5371	-0.484		
+	0.5372	-0.515		
+	0.5373	-0.564		
+	0.5374	-0.54		
+	0.5375	-0.515		
+	0.5376	-0.577		
+	0.5377	-0.446		
+	0.5378	-0.21		
+	0.5379	0.138		
+	0.538	0.68		
+	0.5381	1.756		
+	0.5382	3.043		
+	0.5383	5.015		
+	0.5384	7.764		
+	0.5385	10.993		
+	0.5386	14.489		
+	0.5387	18.382		
+	0.5388	22.855		
+	0.5389	27.47		
+	0.539	32.409		
+	0.5391	37.864		
+	0.5392	43.593		
+	0.5393	49.565		
+	0.5394	55.866		
+	0.5395	62.347		
+	0.5396	68.767		
+	0.5397	75.192		
+	0.5398	81.593		
+	0.5399	87.241		
+	0.54	91.657		
+	0.5401	95.097		
+	0.5402	97.647		
+	0.5403	99.283		
+	0.5404	100.527		
+	0.5405	101.436		
+	0.5406	101.89		
+	0.5407	102.195		
+	0.5408	102.854		
+	0.5409	103.289		
+	0.541	103.974		
+	0.5411	104.72		
+	0.5412	105.516		
+	0.5413	106.219		
+	0.5414	107.009		
+	0.5415	107.874		
+	0.5416	108.508		
+	0.5417	109.037		
+	0.5418	109.721		
+	0.5419	110.001		
+	0.542	110.3		
+	0.5421	110.679		
+	0.5422	110.934		
+	0.5423	111.027		
+	0.5424	111.108		
+	0.5425	111.22		
+	0.5426	111.195		
+	0.5427	111.214		
+	0.5428	111.481		
+	0.5429	111.444		
+	0.543	111.351		
+	0.5431	111.438		
+	0.5432	111.537		
+	0.5433	111.413		
+	0.5434	111.444		
+	0.5435	111.525		
+	0.5436	111.575		
+	0.5437	111.581		
+	0.5438	111.824		
+	0.5439	111.991		
+	0.544	111.923		
+	0.5441	112.147		
+	0.5442	112.24		
+	0.5443	112.159		
+	0.5444	112.01		
+	0.5445	111.805		
+	0.5446	111.295		
+	0.5447	110.287		
+	0.5448	109.093		
+	0.5449	107.202		
+	0.545	104.378		
+	0.5451	100.627		
+	0.5452	95.209		
+	0.5453	86.712		
+	0.5454	77.201		
+	0.5455	69.768		
+	0.5456	63.113		
+	0.5457	56.948		
+	0.5458	51.35		
+	0.5459	46.088		
+	0.546	41.093		
+	0.5461	36.508		
+	0.5462	32.26		
+	0.5463	28.173		
+	0.5464	24.553		
+	0.5465	21.132		
+	0.5466	17.891		
+	0.5467	14.856		
+	0.5468	12.318		
+	0.5469	9.786		
+	0.547	7.441		
+	0.5471	5.513		
+	0.5472	3.759		
+	0.5473	2.16		
+	0.5474	0.866		
+	0.5475	-0.117		
+	0.5476	-1.093		
+	0.5477	-1.852		
+	0.5478	-2.269		
+	0.5479	-2.661		
+	0.548	-2.978		
+	0.5481	-3.152		
+	0.5482	-3.046		
+	0.5483	-3.146		
+	0.5484	-3.165		
+	0.5485	-3.071		
+	0.5486	-2.984		
+	0.5487	-2.966		
+	0.5488	-2.934		
+	0.5489	-2.829		
+	0.549	-2.885		
+	0.5491	-2.804		
+	0.5492	-2.723		
+	0.5493	-2.748		
+	0.5494	-2.686		
+	0.5495	-2.655		
+	0.5496	-2.511		
+	0.5497	-2.543		
+	0.5498	-2.443		
+	0.5499	-2.306		
+	0.55	-2.288		
+	0.5501	-2.238		
+	0.5502	-2.144		
+	0.5503	-2.07		
+	0.5504	-2.12		
+	0.5505	-2.039		
+	0.5506	-1.995		
+	0.5507	-2.051		
+	0.5508	-2.113		
+	0.5509	-1.983		
+	0.551	-1.97		
+	0.5511	-1.952		
+	0.5512	-1.865		
+	0.5513	-1.865		
+	0.5514	-1.84		
+	0.5515	-1.678		
+	0.5516	-1.56		
+	0.5517	-1.56		
+	0.5518	-1.379		
+	0.5519	-1.255		
+	0.552	-1.305		
+	0.5521	-1.205		
+	0.5522	-1.087		
+	0.5523	-1.081		
+	0.5524	-1.112		
+	0.5525	-1.075		
+	0.5526	-1		
+	0.5527	-0.907		
+	0.5528	-0.907		
+	0.5529	-0.813		
+	0.553	-0.77		
+	0.5531	-0.751		
+	0.5532	-0.633		
+	0.5533	-0.564		
+	0.5534	-0.515		
+	0.5535	-0.515		
+	0.5536	-0.465		
+	0.5537	-0.533		
+	0.5538	-0.428		
+	0.5539	-0.316		
+	0.554	-0.086		
+	0.5541	0.132		
+	0.5542	0.742		
+	0.5543	1.494		
+	0.5544	2.72		
+	0.5545	4.536		
+	0.5546	7.23		
+	0.5547	10.253		
+	0.5548	13.736		
+	0.5549	17.667		
+	0.555	21.99		
+	0.5551	26.593		
+	0.5552	31.545		
+	0.5553	36.819		
+	0.5554	42.399		
+	0.5555	48.476		
+	0.5556	54.721		
+	0.5557	61.072		
+	0.5558	67.373		
+	0.5559	73.867		
+	0.556	80.156		
+	0.5561	85.879		
+	0.5562	90.563		
+	0.5563	94.195		
+	0.5564	96.783		
+	0.5565	98.78		
+	0.5566	100.148		
+	0.5567	101.075		
+	0.5568	101.703		
+	0.5569	102.201		
+	0.557	102.748		
+	0.5571	103.215		
+	0.5572	103.83		
+	0.5573	104.633		
+	0.5574	105.274		
+	0.5575	106.057		
+	0.5576	106.847		
+	0.5577	107.612		
+	0.5578	108.166		
+	0.5579	108.869		
+	0.558	109.373		
+	0.5581	109.777		
+	0.5582	110.181		
+	0.5583	110.542		
+	0.5584	110.828		
+	0.5585	110.928		
+	0.5586	111.164		
+	0.5587	111.307		
+	0.5588	111.301		
+	0.5589	111.413		
+	0.559	111.444		
+	0.5591	111.382		
+	0.5592	111.407		
+	0.5593	111.457		
+	0.5594	111.413		
+	0.5595	111.32		
+	0.5596	111.369		
+	0.5597	111.32		
+	0.5598	111.394		
+	0.5599	111.612		
+	0.56	111.743		
+	0.5601	111.886		
+	0.5602	112.023		
+	0.5603	112.215		
+	0.5604	112.315		
+	0.5605	112.321		
+	0.5606	112.315		
+	0.5607	112.023		
+	0.5608	111.5		
+	0.5609	110.741		
+	0.561	109.566		
+	0.5611	107.755		
+	0.5612	105.249		
+	0.5613	101.896		
+	0.5614	96.951		
+	0.5615	89.735		
+	0.5616	80.088		
+	0.5617	72.02		
+	0.5618	65.271		
+	0.5619	59.069		
+	0.562	53.347		
+	0.5621	47.941		
+	0.5622	42.946		
+	0.5623	38.25		
+	0.5624	33.815		
+	0.5625	29.679		
+	0.5626	25.859		
+	0.5627	22.314		
+	0.5628	18.992		
+	0.5629	15.95		
+	0.563	13.164		
+	0.5631	10.632		
+	0.5632	8.256		
+	0.5633	6.247		
+	0.5634	4.48		
+	0.5635	2.732		
+	0.5636	1.426		
+	0.5637	0.4		
+	0.5638	-0.676		
+	0.5639	-1.386		
+	0.564	-1.933		
+	0.5641	-2.493		
+	0.5642	-2.785		
+	0.5643	-3.015		
+	0.5644	-3.084		
+	0.5645	-3.27		
+	0.5646	-3.221		
+	0.5647	-3.152		
+	0.5648	-3.127		
+	0.5649	-3.028		
+	0.565	-2.866		
+	0.5651	-2.841		
+	0.5652	-2.872		
+	0.5653	-2.729		
+	0.5654	-2.648		
+	0.5655	-2.623		
+	0.5656	-2.505		
+	0.5657	-2.48		
+	0.5658	-2.499		
+	0.5659	-2.524		
+	0.566	-2.387		
+	0.5661	-2.375		
+	0.5662	-2.368		
+	0.5663	-2.275		
+	0.5664	-2.163		
+	0.5665	-2.219		
+	0.5666	-2.101		
+	0.5667	-2.008		
+	0.5668	-2.032		
+	0.5669	-2.076		
+	0.567	-1.914		
+	0.5671	-1.896		
+	0.5672	-1.939		
+	0.5673	-1.746		
+	0.5674	-1.809		
+	0.5675	-1.865		
+	0.5676	-1.802		
+	0.5677	-1.634		
+	0.5678	-1.684		
+	0.5679	-1.616		
+	0.568	-1.454		
+	0.5681	-1.41		
+	0.5682	-1.404		
+	0.5683	-1.224		
+	0.5684	-1.143		
+	0.5685	-1.168		
+	0.5686	-1.037		
+	0.5687	-0.863		
+	0.5688	-0.826		
+	0.5689	-0.876		
+	0.569	-0.739		
+	0.5691	-0.708		
+	0.5692	-0.832		
+	0.5693	-0.757		
+	0.5694	-0.639		
+	0.5695	-0.757		
+	0.5696	-0.664		
+	0.5697	-0.577		
+	0.5698	-0.596		
+	0.5699	-0.558		
+	0.57	-0.39		
+	0.5701	-0.322		
+	0.5702	-0.278		
+	0.5703	0.132		
+	0.5704	0.667		
+	0.5705	1.239		
+	0.5706	2.303		
+	0.5707	3.895		
+	0.5708	6.178		
+	0.5709	9.002		
+	0.571	12.311		
+	0.5711	16.044		
+	0.5712	20.074		
+	0.5713	24.541		
+	0.5714	29.374		
+	0.5715	34.449		
+	0.5716	40.029		
+	0.5717	45.926		
+	0.5718	52.034		
+	0.5719	58.298		
+	0.572	64.711		
+	0.5721	71.149		
+	0.5722	77.425		
+	0.5723	83.434		
+	0.5724	88.647		
+	0.5725	92.584		
+	0.5726	95.595		
+	0.5727	97.94		
+	0.5728	99.538		
+	0.5729	100.459		
+	0.573	101.274		
+	0.5731	101.884		
+	0.5732	102.269		
+	0.5733	102.947		
+	0.5734	103.588		
+	0.5735	104.166		
+	0.5736	104.969		
+	0.5737	105.883		
+	0.5738	106.574		
+	0.5739	107.258		
+	0.574	107.998		
+	0.5741	108.707		
+	0.5742	109.13		
+	0.5743	109.547		
+	0.5744	110.113		
+	0.5745	110.312		
+	0.5746	110.53		
+	0.5747	110.872		
+	0.5748	111.052		
+	0.5749	111.108		
+	0.575	111.282		
+	0.5751	111.438		
+	0.5752	111.401		
+	0.5753	111.494		
+	0.5754	111.637		
+	0.5755	111.593		
+	0.5756	111.575		
+	0.5757	111.6		
+	0.5758	111.575		
+	0.5759	111.444		
+	0.576	111.587		
+	0.5761	111.68		
+	0.5762	111.699		
+	0.5763	111.824		
+	0.5764	112.159		
+	0.5765	112.166		
+	0.5766	112.302		
+	0.5767	112.489		
+	0.5768	112.47		
+	0.5769	112.278		
+	0.577	112.085		
+	0.5771	111.606		
+	0.5772	110.505		
+	0.5773	109.012		
+	0.5774	107.077		
+	0.5775	104.061		
+	0.5776	99.986		
+	0.5777	94.481		
+	0.5778	85.636		
+	0.5779	76.374		
+	0.578	69.059		
+	0.5781	62.752		
+	0.5782	56.612		
+	0.5783	51.101		
+	0.5784	45.988		
+	0.5785	41.099		
+	0.5786	36.428		
+	0.5787	32.303		
+	0.5788	28.36		
+	0.5789	24.553		
+	0.579	21.151		
+	0.5791	18.034		
+	0.5792	14.893		
+	0.5793	12.125		
+	0.5794	9.798		
+	0.5795	7.466		
+	0.5796	5.457		
+	0.5797	3.808		
+	0.5798	2.235		
+	0.5799	0.866		
+	0.58	-0.073		
+	0.5801	-0.838		
+	0.5802	-1.622		
+	0.5803	-2.176		
+	0.5804	-2.431		
+	0.5805	-2.729		
+	0.5806	-3.009		
+	0.5807	-2.99		
+	0.5808	-3.059		
+	0.5809	-3.165		
+	0.581	-3.14		
+	0.5811	-2.966		
+	0.5812	-3.034		
+	0.5813	-3.003		
+	0.5814	-2.903		
+	0.5815	-2.866		
+	0.5816	-2.76		
+	0.5817	-2.679		
+	0.5818	-2.493		
+	0.5819	-2.561		
+	0.582	-2.474		
+	0.5821	-2.275		
+	0.5822	-2.356		
+	0.5823	-2.387		
+	0.5824	-2.232		
+	0.5825	-2.225		
+	0.5826	-2.325		
+	0.5827	-2.132		
+	0.5828	-2.132		
+	0.5829	-2.207		
+	0.583	-2.151		
+	0.5831	-2.039		
+	0.5832	-2.051		
+	0.5833	-2.045		
+	0.5834	-1.815		
+	0.5835	-1.815		
+	0.5836	-1.858		
+	0.5837	-1.697		
+	0.5838	-1.634		
+	0.5839	-1.665		
+	0.584	-1.554		
+	0.5841	-1.485		
+	0.5842	-1.473		
+	0.5843	-1.554		
+	0.5844	-1.354		
+	0.5845	-1.292		
+	0.5846	-1.317		
+	0.5847	-1.118		
+	0.5848	-1.087		
+	0.5849	-1.019		
+	0.585	-0.95		
+	0.5851	-0.776		
+	0.5852	-0.82		
+	0.5853	-0.826		
+	0.5854	-0.639		
+	0.5855	-0.552		
+	0.5856	-0.701		
+	0.5857	-0.62		
+	0.5858	-0.502		
+	0.5859	-0.664		
+	0.586	-0.602		
+	0.5861	-0.428		
+	0.5862	-0.49		
+	0.5863	-0.54		
+	0.5864	-0.328		
+	0.5865	-0.129		
+	0.5866	0.219		
+	0.5867	0.922		
+	0.5868	1.868		
+	0.5869	3.012		
+	0.587	4.972		
+	0.5871	7.814		
+	0.5872	10.949		
+	0.5873	14.314		
+	0.5874	18.271		
+	0.5875	22.494		
+	0.5876	26.985		
+	0.5877	32.073		
+	0.5878	37.392		
+	0.5879	42.897		
+	0.588	48.881		
+	0.5881	55.169		
+	0.5882	61.433		
+	0.5883	67.747		
+	0.5884	74.259		
+	0.5885	80.492		
+	0.5886	86.034		
+	0.5887	90.712		
+	0.5888	94.388		
+	0.5889	96.895		
+	0.589	98.761		
+	0.5891	100.167		
+	0.5892	101.013		
+	0.5893	101.597		
+	0.5894	102.157		
+	0.5895	102.686		
+	0.5896	103.096		
+	0.5897	103.762		
+	0.5898	104.62		
+	0.5899	105.342		
+	0.59	106.151		
+	0.5901	107.109		
+	0.5902	107.724		
+	0.5903	108.433		
+	0.5904	109.062		
+	0.5905	109.634		
+	0.5906	109.945		
+	0.5907	110.318		
+	0.5908	110.685		
+	0.5909	110.822		
+	0.591	110.99		
+	0.5911	111.307		
+	0.5912	111.382		
+	0.5913	111.338		
+	0.5914	111.556		
+	0.5915	111.693		
+	0.5916	111.643		
+	0.5917	111.755		
+	0.5918	111.898		
+	0.5919	111.792		
+	0.592	111.824		
+	0.5921	111.935		
+	0.5922	111.96		
+	0.5923	111.911		
+	0.5924	112.029		
+	0.5925	112.147		
+	0.5926	112.178		
+	0.5927	112.377		
+	0.5928	112.62		
+	0.5929	112.626		
+	0.593	112.607		
+	0.5931	112.701		
+	0.5932	112.557		
+	0.5933	111.998		
+	0.5934	111.519		
+	0.5935	110.48		
+	0.5936	108.676		
+	0.5937	106.412		
+	0.5938	103.314		
+	0.5939	98.68		
+	0.594	92.062		
+	0.5941	82.551		
+	0.5942	74.01		
+	0.5943	67.031		
+	0.5944	60.823		
+	0.5945	55.07		
+	0.5946	49.459		
+	0.5947	44.346		
+	0.5948	39.737		
+	0.5949	35.277		
+	0.595	31.115		
+	0.5951	27.383		
+	0.5952	23.726		
+	0.5953	20.249		
+	0.5954	17.188		
+	0.5955	14.445		
+	0.5956	11.665		
+	0.5957	9.12		
+	0.5958	7.136		
+	0.5959	5.115		
+	0.596	3.354		
+	0.5961	1.924		
+	0.5962	0.742		
+	0.5963	-0.421		
+	0.5964	-1.205		
+	0.5965	-1.734		
+	0.5966	-2.238		
+	0.5967	-2.661		
+	0.5968	-2.686		
+	0.5969	-2.903		
+	0.597	-3.084		
+	0.5971	-3.015		
+	0.5972	-2.885		
+	0.5973	-3.015		
+	0.5974	-2.99		
+	0.5975	-2.928		
+	0.5976	-2.953		
+	0.5977	-2.816		
+	0.5978	-2.742		
+	0.5979	-2.791		
+	0.598	-2.698		
+	0.5981	-2.599		
+	0.5982	-2.418		
+	0.5983	-2.468		
+	0.5984	-2.368		
+	0.5985	-2.194		
+	0.5986	-2.244		
+	0.5987	-2.238		
+	0.5988	-2.076		
+	0.5989	-2.126		
+	0.599	-2.107		
+	0.5991	-2.07		
+	0.5992	-1.989		
+	0.5993	-2.151		
+	0.5994	-2.014		
+	0.5995	-1.958		
+	0.5996	-2.001		
+	0.5997	-2.001		
+	0.5998	-1.833		
+	0.5999	-1.74		
+	0.6	-1.74		
+	0.6001	-1.572		
+	0.6002	-1.541		
+	0.6003	-1.554		
+	0.6004	-1.435		
+	0.6005	-1.342		
+	0.6006	-1.267		
+	0.6007	-1.286		
+	0.6008	-1.199		
+	0.6009	-1.099		
+	0.601	-1.193		
+	0.6011	-1.056		
+	0.6012	-0.969		
+	0.6013	-0.981		
+	0.6014	-0.876		
+	0.6015	-0.726		
+	0.6016	-0.701		
+	0.6017	-0.683		
+	0.6018	-0.564		
+	0.6019	-0.515		
+	0.602	-0.54		
+	0.6021	-0.533		
+	0.6022	-0.421		
+	0.6023	-0.434		
+	0.6024	-0.527		
+	0.6025	-0.378		
+	0.6026	-0.334		
+	0.6027	-0.316		
+	0.6028	0.02		
+	0.6029	0.393		
+	0.603	0.991		
+	0.6031	1.936		
+	0.6032	3.553		
+	0.6033	5.587		
+	0.6034	8.424		
+	0.6035	11.665		
+	0.6036	15.21		
+	0.6037	19.154		
+	0.6038	23.545		
+	0.6039	28.229		
+	0.604	33.199		
+	0.6041	38.518		
+	0.6042	44.259		
+	0.6043	50.106		
+	0.6044	56.283		
+	0.6045	62.727		
+	0.6046	68.966		
+	0.6047	75.242		
+	0.6048	81.462		
+	0.6049	87.011		
+	0.605	91.508		
+	0.6051	94.942		
+	0.6052	97.43		
+	0.6053	99.296		
+	0.6054	100.478		
+	0.6055	101.473		
+	0.6056	102.07		
+	0.6057	102.437		
+	0.6058	103.016		
+	0.6059	103.582		
+	0.606	104.092		
+	0.6061	104.844		
+	0.6062	105.697		
+	0.6063	106.468		
+	0.6064	107.245		
+	0.6065	108.017		
+	0.6066	108.794		
+	0.6067	109.304		
+	0.6068	109.883		
+	0.6069	110.356		
+	0.607	110.648		
+	0.6071	110.953		
+	0.6072	111.332		
+	0.6073	111.519		
+	0.6074	111.531		
+	0.6075	111.774		
+	0.6076	111.848		
+	0.6077	111.867		
+	0.6078	111.929		
+	0.6079	112.035		
+	0.608	111.96		
+	0.6081	112.023		
+	0.6082	112.116		
+	0.6083	112.141		
+	0.6084	112.191		
+	0.6085	112.271		
+	0.6086	112.327		
+	0.6087	112.433		
+	0.6088	112.613		
+	0.6089	112.781		
+	0.609	112.875		
+	0.6091	112.999		
+	0.6092	113.161		
+	0.6093	113.18		
+	0.6094	113.08		
+	0.6095	113.012		
+	0.6096	112.533		
+	0.6097	111.861		
+	0.6098	110.803		
+	0.6099	109.143		
+	0.61	106.798		
+	0.6101	103.644		
+	0.6102	99.091		
+	0.6103	92.572		
+	0.6104	83.024		
+	0.6105	74.608		
+	0.6106	67.778		
+	0.6107	61.371		
+	0.6108	55.505		
+	0.6109	50.1		
+	0.611	44.999		
+	0.6111	40.234		
+	0.6112	35.756		
+	0.6113	31.613		
+	0.6114	27.688		
+	0.6115	24.049		
+	0.6116	20.728		
+	0.6117	17.543		
+	0.6118	14.663		
+	0.6119	12.056		
+	0.612	9.618		
+	0.6121	7.354		
+	0.6122	5.475		
+	0.6123	3.696		
+	0.6124	2.185		
+	0.6125	0.991		
+	0.6126	-0.104		
+	0.6127	-1.012		
+	0.6128	-1.709		
+	0.6129	-2.157		
+	0.613	-2.555		
+	0.6131	-2.86		
+	0.6132	-2.941		
+	0.6133	-2.934		
+	0.6134	-3.009		
+	0.6135	-2.978		
+	0.6136	-2.878		
+	0.6137	-2.829		
+	0.6138	-2.866		
+	0.6139	-2.742		
+	0.614	-2.735		
+	0.6141	-2.71		
+	0.6142	-2.642		
+	0.6143	-2.574		
+	0.6144	-2.555		
+	0.6145	-2.474		
+	0.6146	-2.487		
+	0.6147	-2.387		
+	0.6148	-2.393		
+	0.6149	-2.263		
+	0.615	-2.132		
+	0.6151	-2.151		
+	0.6152	-2.107		
+	0.6153	-2.02		
+	0.6154	-2.001		
+	0.6155	-1.958		
+	0.6156	-1.939		
+	0.6157	-1.933		
+	0.6158	-1.989		
+	0.6159	-1.939		
+	0.616	-1.858		
+	0.6161	-1.846		
+	0.6162	-1.74		
+	0.6163	-1.709		
+	0.6164	-1.647		
+	0.6165	-1.597		
+	0.6166	-1.498		
+	0.6167	-1.386		
+	0.6168	-1.342		
+	0.6169	-1.274		
+	0.617	-1.218		
+	0.6171	-1.174		
+	0.6172	-1.087		
+	0.6173	-0.975		
+	0.6174	-0.981		
+	0.6175	-0.931		
+	0.6176	-0.894		
+	0.6177	-0.788		
+	0.6178	-0.732		
+	0.6179	-0.695		
+	0.618	-0.676		
+	0.6181	-0.633		
+	0.6182	-0.533		
+	0.6183	-0.365		
+	0.6184	-0.434		
+	0.6185	-0.434		
+	0.6186	-0.328		
+	0.6187	-0.309		
+	0.6188	-0.272		
+	0.6189	-0.185		
+	0.619	-0.067		
+	0.6191	0.182		
+	0.6192	0.617		
+	0.6193	1.407		
+	0.6194	2.552		
+	0.6195	4.244		
+	0.6196	6.614		
+	0.6197	9.587		
+	0.6198	12.809		
+	0.6199	16.61		
+	0.62	20.765		
+	0.6201	25.194		
+	0.6202	29.94		
+	0.6203	35.103		
+	0.6204	40.508		
+	0.6205	46.243		
+	0.6206	52.333		
+	0.6207	58.59		
+	0.6208	64.736		
+	0.6209	71.006		
+	0.621	77.351		
+	0.6211	83.285		
+	0.6212	88.466		
+	0.6213	92.702		
+	0.6214	95.844		
+	0.6215	98.064		
+	0.6216	99.831		
+	0.6217	101		
+	0.6218	101.734		
+	0.6219	102.362		
+	0.622	102.916		
+	0.6221	103.345		
+	0.6222	103.936		
+	0.6223	104.614		
+	0.6224	105.373		
+	0.6225	106.039		
+	0.6226	106.816		
+	0.6227	107.78		
+	0.6228	108.384		
+	0.6229	109.062		
+	0.623	109.671		
+	0.6231	110.094		
+	0.6232	110.567		
+	0.6233	110.984		
+	0.6234	111.239		
+	0.6235	111.519		
+	0.6236	111.749		
+	0.6237	111.948		
+	0.6238	111.979		
+	0.6239	112.11		
+	0.624	112.191		
+	0.6241	112.191		
+	0.6242	112.271		
+	0.6243	112.296		
+	0.6244	112.365		
+	0.6245	112.346		
+	0.6246	112.278		
+	0.6247	112.421		
+	0.6248	112.396		
+	0.6249	112.489		
+	0.625	112.763		
+	0.6251	112.987		
+	0.6252	113.049		
+	0.6253	113.323		
+	0.6254	113.522		
+	0.6255	113.559		
+	0.6256	113.584		
+	0.6257	113.54		
+	0.6258	113.217		
+	0.6259	112.719		
+	0.626	111.985		
+	0.6261	110.754		
+	0.6262	108.944		
+	0.6263	106.487		
+	0.6264	103.04		
+	0.6265	98.195		
+	0.6266	91.035		
+	0.6267	81.556		
+	0.6268	73.444		
+	0.6269	66.745		
+	0.627	60.631		
+	0.6271	54.852		
+	0.6272	49.44		
+	0.6273	44.458		
+	0.6274	39.78		
+	0.6275	35.351		
+	0.6276	31.178		
+	0.6277	27.47		
+	0.6278	23.775		
+	0.6279	20.398		
+	0.628	17.269		
+	0.6281	14.402		
+	0.6282	11.652		
+	0.6283	9.382		
+	0.6284	7.267		
+	0.6285	5.27		
+	0.6286	3.547		
+	0.6287	2.172		
+	0.6288	0.891		
+	0.6289	-0.16		
+	0.629	-0.913		
+	0.6291	-1.572		
+	0.6292	-2.182		
+	0.6293	-2.499		
+	0.6294	-2.723		
+	0.6295	-2.922		
+	0.6296	-3.04		
+	0.6297	-2.997		
+	0.6298	-3.028		
+	0.6299	-3.015		
+	0.63	-2.86		
+	0.6301	-2.748		
+	0.6302	-2.735		
+	0.6303	-2.717		
+	0.6304	-2.574		
+	0.6305	-2.53		
+	0.6306	-2.561		
+	0.6307	-2.387		
+	0.6308	-2.362		
+	0.6309	-2.443		
+	0.631	-2.325		
+	0.6311	-2.232		
+	0.6312	-2.256		
+	0.6313	-2.194		
+	0.6314	-2.176		
+	0.6315	-2.144		
+	0.6316	-2.101		
+	0.6317	-1.933		
+	0.6318	-1.902		
+	0.6319	-2.014		
+	0.632	-1.84		
+	0.6321	-1.784		
+	0.6322	-1.809		
+	0.6323	-1.79		
+	0.6324	-1.703		
+	0.6325	-1.721		
+	0.6326	-1.759		
+	0.6327	-1.566		
+	0.6328	-1.491		
+	0.6329	-1.547		
+	0.633	-1.448		
+	0.6331	-1.361		
+	0.6332	-1.323		
+	0.6333	-1.149		
+	0.6334	-1		
+	0.6335	-1		
+	0.6336	-0.981		
+	0.6337	-0.813		
+	0.6338	-0.826		
+	0.6339	-0.844		
+	0.634	-0.708		
+	0.6341	-0.589		
+	0.6342	-0.664		
+	0.6343	-0.602		
+	0.6344	-0.44		
+	0.6345	-0.496		
+	0.6346	-0.54		
+	0.6347	-0.459		
+	0.6348	-0.403		
+	0.6349	-0.372		
+	0.635	-0.365		
+	0.6351	-0.197		
+	0.6352	-0.191		
+	0.6353	0.026		
+	0.6354	0.456		
+	0.6355	0.959		
+	0.6356	1.749		
+	0.6357	3.13		
+	0.6358	4.947		
+	0.6359	7.472		
+	0.636	10.545		
+	0.6361	14.122		
+	0.6362	17.798		
+	0.6363	21.965		
+	0.6364	26.637		
+	0.6365	31.433		
+	0.6366	36.558		
+	0.6367	42.169		
+	0.6368	48.109		
+	0.6369	54.037		
+	0.637	60.363		
+	0.6371	66.677		
+	0.6372	72.86		
+	0.6373	78.993		
+	0.6374	84.896		
+	0.6375	89.76		
+	0.6376	93.542		
+	0.6377	96.559		
+	0.6378	98.724		
+	0.6379	100.098		
+	0.638	101.168		
+	0.6381	102.039		
+	0.6382	102.537		
+	0.6383	103.016		
+	0.6384	103.675		
+	0.6385	104.253		
+	0.6386	104.851		
+	0.6387	105.653		
+	0.6388	106.555		
+	0.6389	107.189		
+	0.639	107.998		
+	0.6391	108.813		
+	0.6392	109.373		
+	0.6393	109.858		
+	0.6394	110.48		
+	0.6395	110.822		
+	0.6396	111.058		
+	0.6397	111.338		
+	0.6398	111.736		
+	0.6399	111.811		
+	0.64	112.029		
+	0.6401	112.278		
+	0.6402	112.259		
+	0.6403	112.246		
+	0.6404	112.489		
+	0.6405	112.526		
+	0.6406	112.414		
+	0.6407	112.545		
+	0.6408	112.595		
+	0.6409	112.477		
+	0.641	112.489		
+	0.6411	112.757		
+	0.6412	112.744		
+	0.6413	112.8		
+	0.6414	113.13		
+	0.6415	113.372		
+	0.6416	113.428		
+	0.6417	113.69		
+	0.6418	113.907		
+	0.6419	113.82		
+	0.642	113.714		
+	0.6421	113.547		
+	0.6422	113.005		
+	0.6423	112.159		
+	0.6424	110.872		
+	0.6425	108.962		
+	0.6426	106.175		
+	0.6427	102.742		
+	0.6428	97.716		
+	0.6429	89.853		
+	0.643	80.305		
+	0.6431	72.76		
+	0.6432	66.173		
+	0.6433	59.965		
+	0.6434	54.435		
+	0.6435	49.179		
+	0.6436	44.06		
+	0.6437	39.494		
+	0.6438	35.208		
+	0.6439	31.003		
+	0.644	27.259		
+	0.6441	23.701		
+	0.6442	20.292		
+	0.6443	17.064		
+	0.6444	14.364		
+	0.6445	11.714		
+	0.6446	9.189		
+	0.6447	7.043		
+	0.6448	5.27		
+	0.6449	3.497		
+	0.645	2.011		
+	0.6451	0.953		
+	0.6452	-0.104		
+	0.6453	-1.062		
+	0.6454	-1.566		
+	0.6455	-2.014		
+	0.6456	-2.449		
+	0.6457	-2.698		
+	0.6458	-2.804		
+	0.6459	-2.959		
+	0.646	-3.028		
+	0.6461	-2.922		
+	0.6462	-2.928		
+	0.6463	-2.984		
+	0.6464	-2.822		
+	0.6465	-2.704		
+	0.6466	-2.773		
+	0.6467	-2.623		
+	0.6468	-2.431		
+	0.6469	-2.487		
+	0.647	-2.462		
+	0.6471	-2.263		
+	0.6472	-2.238		
+	0.6473	-2.294		
+	0.6474	-2.163		
+	0.6475	-2.07		
+	0.6476	-2.176		
+	0.6477	-2.132		
+	0.6478	-2.02		
+	0.6479	-1.983		
+	0.648	-2.07		
+	0.6481	-1.958		
+	0.6482	-1.877		
+	0.6483	-1.933		
+	0.6484	-1.777		
+	0.6485	-1.659		
+	0.6486	-1.74		
+	0.6487	-1.665		
+	0.6488	-1.522		
+	0.6489	-1.572		
+	0.649	-1.547		
+	0.6491	-1.448		
+	0.6492	-1.398		
+	0.6493	-1.448		
+	0.6494	-1.28		
+	0.6495	-1.162		
+	0.6496	-1.274		
+	0.6497	-1.174		
+	0.6498	-0.981		
+	0.6499	-0.994		
+	0.65	-0.95		
+	0.6501	-0.714		
+	0.6502	-0.645		
+	0.6503	-0.695		
+	0.6504	-0.558		
+	0.6505	-0.459		
+	0.6506	-0.533		
+	0.6507	-0.509		
+	0.6508	-0.347		
+	0.6509	-0.403		
+	0.651	-0.502		
+	0.6511	-0.334		
+	0.6512	-0.347		
+	0.6513	-0.453		
+	0.6514	-0.303		
+	0.6515	-0.067		
+	0.6516	0.033		
+	0.6517	0.443		
+	0.6518	1.071		
+	0.6519	1.973		
+	0.652	3.255		
+	0.6521	5.301		
+	0.6522	8.032		
+	0.6523	10.974		
+	0.6524	14.408		
+	0.6525	18.37		
+	0.6526	22.469		
+	0.6527	26.998		
+	0.6528	31.968		
+	0.6529	37.155		
+	0.653	42.617		
+	0.6531	48.545		
+	0.6532	54.628		
+	0.6533	60.73		
+	0.6534	67.075		
+	0.6535	73.382		
+	0.6536	79.416		
+	0.6537	85.101		
+	0.6538	90.109		
+	0.6539	93.878		
+	0.654	96.64		
+	0.6541	98.773		
+	0.6542	100.297		
+	0.6543	101.243		
+	0.6544	101.983		
+	0.6545	102.649		
+	0.6546	103.04		
+	0.6547	103.463		
+	0.6548	104.229		
+	0.6549	104.869		
+	0.655	105.622		
+	0.6551	106.524		
+	0.6552	107.32		
+	0.6553	108.004		
+	0.6554	108.732		
+	0.6555	109.478		
+	0.6556	109.976		
+	0.6557	110.399		
+	0.6558	110.816		
+	0.6559	111.17		
+	0.656	111.332		
+	0.6561	111.687		
+	0.6562	111.898		
+	0.6563	111.879		
+	0.6564	112.147		
+	0.6565	112.296		
+	0.6566	112.321		
+	0.6567	112.358		
+	0.6568	112.564		
+	0.6569	112.557		
+	0.657	112.589		
+	0.6571	112.589		
+	0.6572	112.744		
+	0.6573	112.676		
+	0.6574	112.732		
+	0.6575	112.881		
+	0.6576	112.924		
+	0.6577	113.105		
+	0.6578	113.329		
+	0.6579	113.528		
+	0.658	113.584		
+	0.6581	113.77		
+	0.6582	113.851		
+	0.6583	113.814		
+	0.6584	113.515		
+	0.6585	113.136		
+	0.6586	112.253		
+	0.6587	110.915		
+	0.6588	109.18		
+	0.6589	106.592		
+	0.659	102.935		
+	0.6591	98.039		
+	0.6592	90.569		
+	0.6593	80.921		
+	0.6594	73.133		
+	0.6595	66.646		
+	0.6596	60.351		
+	0.6597	54.659		
+	0.6598	49.415		
+	0.6599	44.514		
+	0.66	39.836		
+	0.6601	35.463		
+	0.6602	31.507		
+	0.6603	27.62		
+	0.6604	23.943		
+	0.6605	20.734		
+	0.6606	17.599		
+	0.6607	14.601		
+	0.6608	11.988		
+	0.6609	9.537		
+	0.661	7.236		
+	0.6611	5.345		
+	0.6612	3.709		
+	0.6613	2.172		
+	0.6614	0.848		
+	0.6615	-0.054		
+	0.6616	-0.807		
+	0.6617	-1.572		
+	0.6618	-2.001		
+	0.6619	-2.343		
+	0.662	-2.636		
+	0.6621	-2.841		
+	0.6622	-2.81		
+	0.6623	-2.903		
+	0.6624	-2.966		
+	0.6625	-2.903		
+	0.6626	-2.847		
+	0.6627	-2.878		
+	0.6628	-2.816		
+	0.6629	-2.729		
+	0.663	-2.71		
+	0.6631	-2.667		
+	0.6632	-2.468		
+	0.6633	-2.418		
+	0.6634	-2.418		
+	0.6635	-2.263		
+	0.6636	-2.194		
+	0.6637	-2.2		
+	0.6638	-2.144		
+	0.6639	-2.001		
+	0.664	-2.045		
+	0.6641	-2.039		
+	0.6642	-1.952		
+	0.6643	-1.989		
+	0.6644	-2.008		
+	0.6645	-1.945		
+	0.6646	-1.877		
+	0.6647	-1.902		
+	0.6648	-1.827		
+	0.6649	-1.709		
+	0.665	-1.665		
+	0.6651	-1.609		
+	0.6652	-1.547		
+	0.6653	-1.466		
+	0.6654	-1.504		
+	0.6655	-1.323		
+	0.6656	-1.267		
+	0.6657	-1.249		
+	0.6658	-1.211		
+	0.6659	-1.099		
+	0.666	-1.131		
+	0.6661	-1.081		
+	0.6662	-0.956		
+	0.6663	-0.857		
+	0.6664	-0.851		
+	0.6665	-0.776		
+	0.6666	-0.602		
+	0.6667	-0.627		
+	0.6668	-0.453		
+	0.6669	-0.403		
+	0.667	-0.434		
+	0.6671	-0.403		
+	0.6672	-0.272		
+	0.6673	-0.297		
+	0.6674	-0.39		
+	0.6675	-0.272		
+	0.6676	-0.266		
+	0.6677	-0.272		
+	0.6678	-0.079		
+	0.6679	0.188		
+	0.668	0.536		
+	0.6681	1.165		
+	0.6682	2.235		
+	0.6683	3.715		
+	0.6684	5.836		
+	0.6685	8.778		
+	0.6686	11.907		
+	0.6687	15.403		
+	0.6688	19.316		
+	0.6689	23.738		
+	0.669	28.217		
+	0.6691	33.056		
+	0.6692	38.412		
+	0.6693	43.96		
+	0.6694	49.776		
+	0.6695	55.791		
+	0.6696	62.067		
+	0.6697	68.207		
+	0.6698	74.452		
+	0.6699	80.523		
+	0.67	86.14		
+	0.6701	90.687		
+	0.6702	94.313		
+	0.6703	97.025		
+	0.6704	98.948		
+	0.6705	100.384		
+	0.6706	101.355		
+	0.6707	102.027		
+	0.6708	102.562		
+	0.6709	103.028		
+	0.671	103.613		
+	0.6711	104.166		
+	0.6712	104.894		
+	0.6713	105.603		
+	0.6714	106.406		
+	0.6715	107.158		
+	0.6716	108.042		
+	0.6717	108.776		
+	0.6718	109.404		
+	0.6719	109.982		
+	0.672	110.461		
+	0.6721	110.735		
+	0.6722	111.251		
+	0.6723	111.457		
+	0.6724	111.662		
+	0.6725	111.724		
+	0.6726	111.942		
+	0.6727	112.072		
+	0.6728	112.041		
+	0.6729	112.222		
+	0.673	112.284		
+	0.6731	112.24		
+	0.6732	112.302		
+	0.6733	112.464		
+	0.6734	112.495		
+	0.6735	112.57		
+	0.6736	112.651		
+	0.6737	112.757		
+	0.6738	112.875		
+	0.6739	112.993		
+	0.674	113.161		
+	0.6741	113.323		
+	0.6742	113.422		
+	0.6743	113.665		
+	0.6744	113.708		
+	0.6745	113.64		
+	0.6746	113.596		
+	0.6747	113.329		
+	0.6748	112.701		
+	0.6749	111.923		
+	0.675	110.573		
+	0.6751	108.57		
+	0.6752	105.877		
+	0.6753	102.163		
+	0.6754	96.969		
+	0.6755	88.852		
+	0.6756	79.64		
+	0.6757	72.138		
+	0.6758	65.482		
+	0.6759	59.467		
+	0.676	53.944		
+	0.6761	48.681		
+	0.6762	43.687		
+	0.6763	39.146		
+	0.6764	34.848		
+	0.6765	30.823		
+	0.6766	27.103		
+	0.6767	23.589		
+	0.6768	20.224		
+	0.6769	17.163		
+	0.677	14.333		
+	0.6771	11.646		
+	0.6772	9.301		
+	0.6773	7.223		
+	0.6774	5.202		
+	0.6775	3.454		
+	0.6776	2.073		
+	0.6777	0.885		
+	0.6778	-0.173		
+	0.6779	-1.031		
+	0.678	-1.572		
+	0.6781	-2.107		
+	0.6782	-2.474		
+	0.6783	-2.605		
+	0.6784	-2.779		
+	0.6785	-2.86		
+	0.6786	-2.891		
+	0.6787	-2.86		
+	0.6788	-2.847		
+	0.6789	-2.829		
+	0.679	-2.692		
+	0.6791	-2.698		
+	0.6792	-2.704		
+	0.6793	-2.567		
+	0.6794	-2.611		
+	0.6795	-2.567		
+	0.6796	-2.412		
+	0.6797	-2.368		
+	0.6798	-2.387		
+	0.6799	-2.281		
+	0.68	-2.169		
+	0.6801	-2.113		
+	0.6802	-2.082		
+	0.6803	-1.989		
+	0.6804	-1.952		
+	0.6805	-1.976		
+	0.6806	-1.952		
+	0.6807	-1.84		
+	0.6808	-1.927		
+	0.6809	-1.858		
+	0.681	-1.809		
+	0.6811	-1.858		
+	0.6812	-1.846		
+	0.6813	-1.759		
+	0.6814	-1.653		
+	0.6815	-1.609		
+	0.6816	-1.504		
+	0.6817	-1.392		
+	0.6818	-1.386		
+	0.6819	-1.305		
+	0.682	-1.162		
+	0.6821	-1.131		
+	0.6822	-1.112		
+	0.6823	-0.981		
+	0.6824	-0.9		
+	0.6825	-0.975		
+	0.6826	-0.869		
+	0.6827	-0.751		
+	0.6828	-0.764		
+	0.6829	-0.72		
+	0.683	-0.54		
+	0.6831	-0.509		
+	0.6832	-0.533		
+	0.6833	-0.378		
+	0.6834	-0.291		
+	0.6835	-0.266		
+	0.6836	-0.26		
+	0.6837	-0.222		
+	0.6838	-0.26		
+	0.6839	-0.229		
+	0.684	-0.123		
+	0.6841	-0.042		
+	0.6842	0.039		
+	0.6843	0.53		
+	0.6844	1.215		
+	0.6845	1.961		
+	0.6846	3.429		
+	0.6847	5.674		
+	0.6848	8.331		
+	0.6849	11.497		
+	0.685	15.092		
+	0.6851	18.967		
+	0.6852	23.066		
+	0.6853	27.694		
+	0.6854	32.664		
+	0.6855	37.796		
+	0.6856	43.239		
+	0.6857	49.123		
+	0.6858	55.032		
+	0.6859	61.147		
+	0.686	67.448		
+	0.6861	73.637		
+	0.6862	79.546		
+	0.6863	85.232		
+	0.6864	90.021		
+	0.6865	93.642		
+	0.6866	96.497		
+	0.6867	98.587		
+	0.6868	100.073		
+	0.6869	101.044		
+	0.687	101.809		
+	0.6871	102.394		
+	0.6872	102.823		
+	0.6873	103.389		
+	0.6874	104.036		
+	0.6875	104.571		
+	0.6876	105.33		
+	0.6877	106.225		
+	0.6878	106.965		
+	0.6879	107.668		
+	0.688	108.433		
+	0.6881	109.13		
+	0.6882	109.615		
+	0.6883	110.113		
+	0.6884	110.691		
+	0.6885	110.984		
+	0.6886	111.195		
+	0.6887	111.556		
+	0.6888	111.718		
+	0.6889	111.724		
+	0.689	112.004		
+	0.6891	112.06		
+	0.6892	112.004		
+	0.6893	112.11		
+	0.6894	112.271		
+	0.6895	112.209		
+	0.6896	112.184		
+	0.6897	112.315		
+	0.6898	112.377		
+	0.6899	112.377		
+	0.69	112.551		
+	0.6901	112.769		
+	0.6902	112.806		
+	0.6903	112.962		
+	0.6904	113.229		
+	0.6905	113.36		
+	0.6906	113.441		
+	0.6907	113.634		
+	0.6908	113.615		
+	0.6909	113.416		
+	0.691	113.242		
+	0.6911	112.8		
+	0.6912	111.867		
+	0.6913	110.598		
+	0.6914	108.807		
+	0.6915	106.219		
+	0.6916	102.773		
+	0.6917	98.07		
+	0.6918	90.625		
+	0.6919	81.095		
+	0.692	73.42		
+	0.6921	66.913		
+	0.6922	60.674		
+	0.6923	54.995		
+	0.6924	49.807		
+	0.6925	44.707		
+	0.6926	39.936		
+	0.6927	35.781		
+	0.6928	31.688		
+	0.6929	27.713		
+	0.693	24.186		
+	0.6931	20.883		
+	0.6932	17.673		
+	0.6933	14.75		
+	0.6934	12.28		
+	0.6935	9.823		
+	0.6936	7.516		
+	0.6937	5.643		
+	0.6938	3.958		
+	0.6939	2.347		
+	0.694	1.165		
+	0.6941	0.089		
+	0.6942	-0.857		
+	0.6943	-1.572		
+	0.6944	-1.908		
+	0.6945	-2.399		
+	0.6946	-2.717		
+	0.6947	-2.773		
+	0.6948	-2.903		
+	0.6949	-2.959		
+	0.695	-2.847		
+	0.6951	-2.816		
+	0.6952	-2.872		
+	0.6953	-2.791		
+	0.6954	-2.611		
+	0.6955	-2.592		
+	0.6956	-2.673		
+	0.6957	-2.524		
+	0.6958	-2.474		
+	0.6959	-2.48		
+	0.696	-2.437		
+	0.6961	-2.337		
+	0.6962	-2.3		
+	0.6963	-2.281		
+	0.6964	-2.144		
+	0.6965	-2.144		
+	0.6966	-2.194		
+	0.6967	-1.958		
+	0.6968	-1.889		
+	0.6969	-1.976		
+	0.697	-1.939		
+	0.6971	-1.734		
+	0.6972	-1.802		
+	0.6973	-1.889		
+	0.6974	-1.709		
+	0.6975	-1.74		
+	0.6976	-1.821		
+	0.6977	-1.634		
+	0.6978	-1.541		
+	0.6979	-1.591		
+	0.698	-1.529		
+	0.6981	-1.404		
+	0.6982	-1.361		
+	0.6983	-1.342		
+	0.6984	-1.131		
+	0.6985	-0.981		
+	0.6986	-1.118		
+	0.6987	-0.919		
+	0.6988	-0.807		
+	0.6989	-0.832		
+	0.699	-0.739		
+	0.6991	-0.602		
+	0.6992	-0.614		
+	0.6993	-0.664		
+	0.6994	-0.477		
+	0.6995	-0.471		
+	0.6996	-0.583		
+	0.6997	-0.434		
+	0.6998	-0.409		
+	0.6999	-0.378		
+	0.7	-0.334		
+	0.7001	-0.135		
+	0.7002	-0.197		
+	0.7003	-0.266		
+	0.7004	0.014		
+	0.7005	0.306		
+	0.7006	0.555		
+	0.7007	1.302		
+	0.7008	2.303		
+	0.7009	3.609		
+	0.701	5.83		
+	0.7011	8.642		
+	0.7012	11.745		
+	0.7013	15.167		
+	0.7014	19.191		
+	0.7015	23.421		
+	0.7016	27.831		
+	0.7017	32.863		
+	0.7018	38.163		
+	0.7019	43.512		
+	0.702	49.31		
+	0.7021	55.374		
+	0.7022	61.439		
+	0.7023	67.485		
+	0.7024	73.637		
+	0.7025	79.646		
+	0.7026	85.139		
+	0.7027	89.909		
+	0.7028	93.654		
+	0.7029	96.279		
+	0.703	98.251		
+	0.7031	99.8		
+	0.7032	100.832		
+	0.7033	101.492		
+	0.7034	102.207		
+	0.7035	102.792		
+	0.7036	103.152		
+	0.7037	103.812		
+	0.7038	104.589		
+	0.7039	105.174		
+	0.704	105.976		
+	0.7041	106.841		
+	0.7042	107.625		
+	0.7043	108.166		
+	0.7044	108.9		
+	0.7045	109.547		
+	0.7046	109.883		
+	0.7047	110.505		
+	0.7048	110.735		
+	0.7049	110.971		
+	0.705	111.208		
+	0.7051	111.544		
+	0.7052	111.693		
+	0.7053	111.705		
+	0.7054	111.911		
+	0.7055	111.991		
+	0.7056	111.942		
+	0.7057	111.991		
+	0.7058	112.147		
+	0.7059	112.091		
+	0.706	112.066		
+	0.7061	112.246		
+	0.7062	112.184		
+	0.7063	112.191		
+	0.7064	112.701		
+	0.7065	112.663		
+	0.7066	112.669		
+	0.7067	112.9		
+	0.7068	113.198		
+	0.7069	113.291		
+	0.707	113.279		
+	0.7071	113.459		
+	0.7072	113.347		
+	0.7073	113.03		
+	0.7074	112.495		
+	0.7075	111.68		
+	0.7076	110.287		
+	0.7077	108.44		
+	0.7078	105.964		
+	0.7079	102.356		
+	0.708	97.361		
+	0.7081	89.878		
+	0.7082	80.647		
+	0.7083	72.841		
+	0.7084	66.428		
+	0.7085	60.419		
+	0.7086	54.703		
+	0.7087	49.409		
+	0.7088	44.676		
+	0.7089	39.892		
+	0.709	35.482		
+	0.7091	31.538		
+	0.7092	27.719		
+	0.7093	23.975		
+	0.7094	20.721		
+	0.7095	17.698		
+	0.7096	14.657		
+	0.7097	11.982		
+	0.7098	9.668		
+	0.7099	7.491		
+	0.71	5.494		
+	0.7101	3.877		
+	0.7102	2.434		
+	0.7103	1.047		
+	0.7104	0.064		
+	0.7105	-0.695		
+	0.7106	-1.466		
+	0.7107	-2.02		
+	0.7108	-2.312		
+	0.7109	-2.636		
+	0.711	-2.928		
+	0.7111	-2.841		
+	0.7112	-2.891		
+	0.7113	-2.99		
+	0.7114	-2.953		
+	0.7115	-2.829		
+	0.7116	-2.847		
+	0.7117	-2.729		
+	0.7118	-2.543		
+	0.7119	-2.586		
+	0.712	-2.524		
+	0.7121	-2.424		
+	0.7122	-2.35		
+	0.7123	-2.356		
+	0.7124	-2.356		
+	0.7125	-2.25		
+	0.7126	-2.306		
+	0.7127	-2.219		
+	0.7128	-2.138		
+	0.7129	-2.088		
+	0.713	-2.101		
+	0.7131	-2.045		
+	0.7132	-1.896		
+	0.7133	-1.939		
+	0.7134	-1.852		
+	0.7135	-1.79		
+	0.7136	-1.802		
+	0.7137	-1.846		
+	0.7138	-1.609		
+	0.7139	-1.653		
+	0.714	-1.672		
+	0.7141	-1.634		
+	0.7142	-1.554		
+	0.7143	-1.578		
+	0.7144	-1.442		
+	0.7145	-1.311		
+	0.7146	-1.342		
+	0.7147	-1.348		
+	0.7148	-1.149		
+	0.7149	-1.025		
+	0.715	-1.006		
+	0.7151	-0.844		
+	0.7152	-0.77		
+	0.7153	-0.751		
+	0.7154	-0.664		
+	0.7155	-0.459		
+	0.7156	-0.502		
+	0.7157	-0.527		
+	0.7158	-0.409		
+	0.7159	-0.428		
+	0.716	-0.459		
+	0.7161	-0.397		
+	0.7162	-0.328		
+	0.7163	-0.365		
+	0.7164	-0.372		
+	0.7165	-0.173		
+	0.7166	-0.185		
+	0.7167	-0.067		
+	0.7168	0.194		
+	0.7169	0.574		
+	0.717	1.115		
+	0.7171	2.073		
+	0.7172	3.528		
+	0.7173	5.556		
+	0.7174	8.144		
+	0.7175	11.291		
+	0.7176	14.632		
+	0.7177	18.37		
+	0.7178	22.618		
+	0.7179	27.134		
+	0.718	31.837		
+	0.7181	37.018		
+	0.7182	42.511		
+	0.7183	48.234		
+	0.7184	54.099		
+	0.7185	60.332		
+	0.7186	66.328		
+	0.7187	72.343		
+	0.7188	78.421		
+	0.7189	84.087		
+	0.719	88.883		
+	0.7191	92.733		
+	0.7192	95.657		
+	0.7193	97.716		
+	0.7194	99.29		
+	0.7195	100.447		
+	0.7196	101.224		
+	0.7197	101.734		
+	0.7198	102.375		
+	0.7199	102.966		
+	0.72	103.463		
+	0.7201	104.173		
+	0.7202	104.919		
+	0.7203	105.74		
+	0.7204	106.487		
+	0.7205	107.376		
+	0.7206	108.085		
+	0.7207	108.626		
+	0.7208	109.205		
+	0.7209	109.74		
+	0.721	110.082		
+	0.7211	110.492		
+	0.7212	110.81		
+	0.7213	111.009		
+	0.7214	111.139		
+	0.7215	111.394		
+	0.7216	111.562		
+	0.7217	111.693		
+	0.7218	111.774		
+	0.7219	111.879		
+	0.722	111.96		
+	0.7221	111.929		
+	0.7222	112.041		
+	0.7223	112.06		
+	0.7224	111.985		
+	0.7225	112.091		
+	0.7226	112.103		
+	0.7227	112.228		
+	0.7228	112.358		
+	0.7229	112.595		
+	0.723	112.669		
+	0.7231	112.837		
+	0.7232	113.03		
+	0.7233	113.242		
+	0.7234	113.211		
+	0.7235	113.167		
+	0.7236	113.018		
+	0.7237	112.539		
+	0.7238	111.824		
+	0.7239	110.673		
+	0.724	108.863		
+	0.7241	106.449		
+	0.7242	103.296		
+	0.7243	98.599		
+	0.7244	91.85		
+	0.7245	82.551		
+	0.7246	74.458		
+	0.7247	67.628		
+	0.7248	61.62		
+	0.7249	55.959		
+	0.725	50.697		
+	0.7251	45.665		
+	0.7252	40.925		
+	0.7253	36.62		
+	0.7254	32.484		
+	0.7255	28.59		
+	0.7256	25.063		
+	0.7257	21.598		
+	0.7258	18.37		
+	0.7259	15.496		
+	0.726	12.691		
+	0.7261	10.215		
+	0.7262	8.044		
+	0.7263	5.998		
+	0.7264	4.2		
+	0.7265	2.639		
+	0.7266	1.42		
+	0.7267	0.356		
+	0.7268	-0.577		
+	0.7269	-1.236		
+	0.727	-1.765		
+	0.7271	-2.232		
+	0.7272	-2.399		
+	0.7273	-2.673		
+	0.7274	-2.81		
+	0.7275	-2.928		
+	0.7276	-2.903		
+	0.7277	-2.86		
+	0.7278	-2.922		
+	0.7279	-2.76		
+	0.728	-2.773		
+	0.7281	-2.748		
+	0.7282	-2.667		
+	0.7283	-2.449		
+	0.7284	-2.455		
+	0.7285	-2.381		
+	0.7286	-2.306		
+	0.7287	-2.25		
+	0.7288	-2.219		
+	0.7289	-2.169		
+	0.729	-2.101		
+	0.7291	-2.107		
+	0.7292	-2.101		
+	0.7293	-2.07		
+	0.7294	-2.032		
+	0.7295	-2.008		
+	0.7296	-1.939		
+	0.7297	-1.989		
+	0.7298	-1.952		
+	0.7299	-1.79		
+	0.73	-1.709		
+	0.7301	-1.715		
+	0.7302	-1.672		
+	0.7303	-1.522		
+	0.7304	-1.547		
+	0.7305	-1.529		
+	0.7306	-1.392		
+	0.7307	-1.392		
+	0.7308	-1.379		
+	0.7309	-1.255		
+	0.731	-1.224		
+	0.7311	-1.168		
+	0.7312	-1.081		
+	0.7313	-1.012		
+	0.7314	-0.913		
+	0.7315	-0.888		
+	0.7316	-0.726		
+	0.7317	-0.627		
+	0.7318	-0.558		
+	0.7319	-0.44		
+	0.732	-0.365		
+	0.7321	-0.397		
+	0.7322	-0.229		
+	0.7323	-0.185		
+	0.7324	-0.21		
+	0.7325	-0.322		
+	0.7326	-0.316		
+	0.7327	-0.241		
+	0.7328	-0.278		
+	0.7329	-0.123		
+	0.733	-0.16		
+	0.7331	0.07		
+	0.7332	0.344		
+	0.7333	1.003		
+	0.7334	1.743		
+	0.7335	3.068		
+	0.7336	4.828		
+	0.7337	7.397		
+	0.7338	10.277		
+	0.7339	13.593		
+	0.734	17.306		
+	0.7341	21.3		
+	0.7342	25.66		
+	0.7343	30.276		
+	0.7344	35.271		
+	0.7345	40.539		
+	0.7346	46.137		
+	0.7347	51.972		
+	0.7348	57.999		
+	0.7349	64.07		
+	0.735	70.26		
+	0.7351	76.212		
+	0.7352	81.96		
+	0.7353	87.185		
+	0.7354	91.409		
+	0.7355	94.606		
+	0.7356	97.044		
+	0.7357	98.748		
+	0.7358	99.993		
+	0.7359	100.832		
+	0.736	101.517		
+	0.7361	102.045		
+	0.7362	102.512		
+	0.7363	103.208		
+	0.7364	103.774		
+	0.7365	104.44		
+	0.7366	105.305		
+	0.7367	106.175		
+	0.7368	106.959		
+	0.7369	107.662		
+	0.737	108.39		
+	0.7371	108.999		
+	0.7372	109.609		
+	0.7373	110.057		
+	0.7374	110.38		
+	0.7375	110.617		
+	0.7376	110.928		
+	0.7377	111.214		
+	0.7378	111.301		
+	0.7379	111.481		
+	0.738	111.562		
+	0.7381	111.643		
+	0.7382	111.662		
+	0.7383	111.892		
+	0.7384	111.935		
+	0.7385	111.873		
+	0.7386	111.998		
+	0.7387	112.091		
+	0.7388	112.079		
+	0.7389	112.141		
+	0.739	112.271		
+	0.7391	112.383		
+	0.7392	112.408		
+	0.7393	112.645		
+	0.7394	112.831		
+	0.7395	112.949		
+	0.7396	113.092		
+	0.7397	113.167		
+	0.7398	113.148		
+	0.7399	113.018		
+	0.74	112.757		
+	0.7401	112.166		
+	0.7402	111.096		
+	0.7403	109.628		
+	0.7404	107.569		
+	0.7405	104.571		
+	0.7406	100.621		
+	0.7407	95.041		
+	0.7408	86.215		
+	0.7409	77.369		
+	0.741	70.372		
+	0.7411	64.126		
+	0.7412	58.149		
+	0.7413	52.718		
+	0.7414	47.699		
+	0.7415	42.729		
+	0.7416	38.374		
+	0.7417	34.244		
+	0.7418	30.232		
+	0.7419	26.531		
+	0.742	23.023		
+	0.7421	19.801		
+	0.7422	16.778		
+	0.7423	13.985		
+	0.7424	11.403		
+	0.7425	8.946		
+	0.7426	6.875		
+	0.7427	5.04		
+	0.7428	3.379		
+	0.7429	1.861		
+	0.743	0.76		
+	0.7431	-0.222		
+	0.7432	-1.099		
+	0.7433	-1.578		
+	0.7434	-1.989		
+	0.7435	-2.319		
+	0.7436	-2.605		
+	0.7437	-2.648		
+	0.7438	-2.723		
+	0.7439	-2.86		
+	0.744	-2.785		
+	0.7441	-2.723		
+	0.7442	-2.829		
+	0.7443	-2.773		
+	0.7444	-2.623		
+	0.7445	-2.679		
+	0.7446	-2.679		
+	0.7447	-2.511		
+	0.7448	-2.505		
+	0.7449	-2.449		
+	0.745	-2.275		
+	0.7451	-2.157		
+	0.7452	-2.275		
+	0.7453	-2.138		
+	0.7454	-2.045		
+	0.7455	-2.008		
+	0.7456	-2.001		
+	0.7457	-1.896		
+	0.7458	-1.952		
+	0.7459	-1.958		
+	0.746	-1.858		
+	0.7461	-1.846		
+	0.7462	-1.883		
+	0.7463	-1.896		
+	0.7464	-1.709		
+	0.7465	-1.753		
+	0.7466	-1.684		
+	0.7467	-1.522		
+	0.7468	-1.435		
+	0.7469	-1.541		
+	0.747	-1.317		
+	0.7471	-1.187		
+	0.7472	-1.249		
+	0.7473	-1.23		
+	0.7474	-1.037		
+	0.7475	-1.081		
+	0.7476	-1.05		
+	0.7477	-0.9		
+	0.7478	-0.813		
+	0.7479	-0.882		
+	0.748	-0.714		
+	0.7481	-0.664		
+	0.7482	-0.639		
+	0.7483	-0.49		
+	0.7484	-0.353		
+	0.7485	-0.297		
+	0.7486	-0.365		
+	0.7487	-0.235		
+	0.7488	-0.173		
+	0.7489	-0.179		
+	0.749	-0.191		
+	0.7491	-0.098		
+	0.7492	-0.266		
+	0.7493	-0.166		
+	0.7494	0.101		
+	0.7495	0.263		
+	0.7496	0.624		
+	0.7497	1.382		
+	0.7498	2.471		
+	0.7499	4.001		
+	0.75	6.352		
+	0.7501	9.195		
+	0.7502	12.243		
+	0.7503	15.776		
+	0.7504	19.832		
+	0.7505	24.024		
+	0.7506	28.385		
+	0.7507	33.348		
+	0.7508	38.511		
+	0.7509	43.805		
+	0.751	49.621		
+	0.7511	55.592		
+	0.7512	61.526		
+	0.7513	67.492		
+	0.7514	73.569		
+	0.7515	79.422		
+	0.7516	84.883		
+	0.7517	89.592		
+	0.7518	93.312		
+	0.7519	95.831		
+	0.752	98.039		
+	0.7521	99.514		
+	0.7522	100.49		
+	0.7523	101.187		
+	0.7524	101.877		
+	0.7525	102.319		
+	0.7526	102.798		
+	0.7527	103.482		
+	0.7528	104.173		
+	0.7529	104.819		
+	0.753	105.578		
+	0.7531	106.487		
+	0.7532	107.283		
+	0.7533	107.973		
+	0.7534	108.8		
+	0.7535	109.366		
+	0.7536	109.69		
+	0.7537	110.206		
+	0.7538	110.617		
+	0.7539	110.778		
+	0.754	111.09		
+	0.7541	111.295		
+	0.7542	111.313		
+	0.7543	111.413		
+	0.7544	111.631		
+	0.7545	111.674		
+	0.7546	111.687		
+	0.7547	111.755		
+	0.7548	111.855		
+	0.7549	111.886		
+	0.755	111.948		
+	0.7551	112.228		
+	0.7552	112.122		
+	0.7553	112.116		
+	0.7554	112.377		
+	0.7555	112.464		
+	0.7556	112.483		
+	0.7557	112.744		
+	0.7558	113.012		
+	0.7559	112.993		
+	0.756	113.099		
+	0.7561	113.304		
+	0.7562	113.005		
+	0.7563	112.75		
+	0.7564	112.365		
+	0.7565	111.587		
+	0.7566	110.287		
+	0.7567	108.539		
+	0.7568	106.126		
+	0.7569	102.611		
+	0.757	97.89		
+	0.7571	90.799		
+	0.7572	81.425		
+	0.7573	73.581		
+	0.7574	67.125		
+	0.7575	61.085		
+	0.7576	55.331		
+	0.7577	50.087		
+	0.7578	45.223		
+	0.7579	40.452		
+	0.758	36.079		
+	0.7581	32.204		
+	0.7582	28.391		
+	0.7583	24.764		
+	0.7584	21.505		
+	0.7585	18.358		
+	0.7586	15.297		
+	0.7587	12.672		
+	0.7588	10.246		
+	0.7589	7.976		
+	0.759	5.948		
+	0.7591	4.262		
+	0.7592	2.627		
+	0.7593	1.239		
+	0.7594	0.325		
+	0.7595	-0.583		
+	0.7596	-1.423		
+	0.7597	-1.933		
+	0.7598	-2.244		
+	0.7599	-2.511		
+	0.76	-2.735		
+	0.7601	-2.679		
+	0.7602	-2.804		
+	0.7603	-2.835		
+	0.7604	-2.791		
+	0.7605	-2.611		
+	0.7606	-2.76		
+	0.7607	-2.661		
+	0.7608	-2.493		
+	0.7609	-2.623		
+	0.761	-2.642		
+	0.7611	-2.449		
+	0.7612	-2.406		
+	0.7613	-2.443		
+	0.7614	-2.281		
+	0.7615	-2.25		
+	0.7616	-2.194		
+	0.7617	-2.188		
+	0.7618	-1.933		
+	0.7619	-1.983		
+	0.762	-1.97		
+	0.7621	-1.771		
+	0.7622	-1.777		
+	0.7623	-1.889		
+	0.7624	-1.84		
+	0.7625	-1.777		
+	0.7626	-1.902		
+	0.7627	-1.796		
+	0.7628	-1.665		
+	0.7629	-1.678		
+	0.763	-1.753		
+	0.7631	-1.522		
+	0.7632	-1.417		
+	0.7633	-1.46		
+	0.7634	-1.249		
+	0.7635	-1.193		
+	0.7636	-1.211		
+	0.7637	-1.155		
+	0.7638	-0.925		
+	0.7639	-0.944		
+	0.764	-0.919		
+	0.7641	-0.857		
+	0.7642	-0.82		
+	0.7643	-0.757		
+	0.7644	-0.714		
+	0.7645	-0.552		
+	0.7646	-0.54		
+	0.7647	-0.577		
+	0.7648	-0.353		
+	0.7649	-0.285		
+	0.765	-0.334		
+	0.7651	-0.129		
+	0.7652	-0.191		
+	0.7653	-0.166		
+	0.7654	-0.123		
+	0.7655	-0.061		
+	0.7656	-0.03		
+	0.7657	-0.017		
+	0.7658	0.281		
+	0.7659	0.487		
+	0.766	1.04		
+	0.7661	2.017		
+	0.7662	3.385		
+	0.7663	5.258		
+	0.7664	8.032		
+	0.7665	11.061		
+	0.7666	14.364		
+	0.7667	18.127		
+	0.7668	22.401		
+	0.7669	26.668		
+	0.767	31.333		
+	0.7671	36.428		
+	0.7672	41.802		
+	0.7673	47.282		
+	0.7674	53.092		
+	0.7675	59.044		
+	0.7676	64.979		
+	0.7677	70.962		
+	0.7678	76.915		
+	0.7679	82.495		
+	0.768	87.477		
+	0.7681	91.676		
+	0.7682	94.823		
+	0.7683	96.945		
+	0.7684	98.761		
+	0.7685	100.16		
+	0.7686	100.894		
+	0.7687	101.56		
+	0.7688	102.188		
+	0.7689	102.611		
+	0.769	103.152		
+	0.7691	103.806		
+	0.7692	104.508		
+	0.7693	105.162		
+	0.7694	106.02		
+	0.7695	106.897		
+	0.7696	107.55		
+	0.7697	108.16		
+	0.7698	108.981		
+	0.7699	109.553		
+	0.77	109.933		
+	0.7701	110.405		
+	0.7702	110.729		
+	0.7703	110.866		
+	0.7704	111.17		
+	0.7705	111.469		
+	0.7706	111.525		
+	0.7707	111.593		
+	0.7708	111.724		
+	0.7709	111.78		
+	0.771	111.712		
+	0.7711	111.867		
+	0.7712	111.904		
+	0.7713	111.836		
+	0.7714	111.892		
+	0.7715	112.147		
+	0.7716	112.172		
+	0.7717	112.234		
+	0.7718	112.52		
+	0.7719	112.595		
+	0.772	112.676		
+	0.7721	112.974		
+	0.7722	113.186		
+	0.7723	113.242		
+	0.7724	113.18		
+	0.7725	113.242		
+	0.7726	113.024		
+	0.7727	112.582		
+	0.7728	111.991		
+	0.7729	110.94		
+	0.773	109.279		
+	0.7731	107.245		
+	0.7732	104.428		
+	0.7733	100.285		
+	0.7734	94.668		
+	0.7735	85.953		
+	0.7736	77.282		
+	0.7737	70.297		
+	0.7738	64.083		
+	0.7739	58.298		
+	0.774	52.824		
+	0.7741	47.724		
+	0.7742	43.002		
+	0.7743	38.374		
+	0.7744	34.232		
+	0.7745	30.332		
+	0.7746	26.562		
+	0.7747	23.004		
+	0.7748	19.913		
+	0.7749	16.902		
+	0.775	14.041		
+	0.7751	11.528		
+	0.7752	9.27		
+	0.7753	7.062		
+	0.7754	5.177		
+	0.7755	3.628		
+	0.7756	2.135		
+	0.7757	0.854		
+	0.7758	-0.104		
+	0.7759	-0.9		
+	0.776	-1.659		
+	0.7761	-2.076		
+	0.7762	-2.3		
+	0.7763	-2.686		
+	0.7764	-2.866		
+	0.7765	-2.847		
+	0.7766	-2.86		
+	0.7767	-2.86		
+	0.7768	-2.773		
+	0.7769	-2.673		
+	0.777	-2.679		
+	0.7771	-2.648		
+	0.7772	-2.511		
+	0.7773	-2.549		
+	0.7774	-2.543		
+	0.7775	-2.418		
+	0.7776	-2.325		
+	0.7777	-2.343		
+	0.7778	-2.281		
+	0.7779	-2.263		
+	0.778	-2.256		
+	0.7781	-2.238		
+	0.7782	-2.051		
+	0.7783	-1.976		
+	0.7784	-1.945		
+	0.7785	-1.796		
+	0.7786	-1.784		
+	0.7787	-1.821		
+	0.7788	-1.74		
+	0.7789	-1.709		
+	0.779	-1.784		
+	0.7791	-1.746		
+	0.7792	-1.628		
+	0.7793	-1.703		
+	0.7794	-1.659		
+	0.7795	-1.504		
+	0.7796	-1.417		
+	0.7797	-1.491		
+	0.7798	-1.373		
+	0.7799	-1.249		
+	0.78	-1.211		
+	0.7801	-1.062		
+	0.7802	-0.931		
+	0.7803	-0.801		
+	0.7804	-0.782		
+	0.7805	-0.652		
+	0.7806	-0.571		
+	0.7807	-0.596		
+	0.7808	-0.577		
+	0.7809	-0.471		
+	0.781	-0.477		
+	0.7811	-0.465		
+	0.7812	-0.353		
+	0.7813	-0.285		
+	0.7814	-0.403		
+	0.7815	-0.154		
+	0.7816	-0.179		
+	0.7817	-0.129		
+	0.7818	-0.104		
+	0.7819	0.008		
+	0.782	0.051		
+	0.7821	0.163		
+	0.7822	0.574		
+	0.7823	0.922		
+	0.7824	1.588		
+	0.7825	2.745		
+	0.7826	4.449		
+	0.7827	6.813		
+	0.7828	9.649		
+	0.7829	12.853		
+	0.783	16.404		
+	0.7831	20.298		
+	0.7832	24.696		
+	0.7833	29.224		
+	0.7834	34.089		
+	0.7835	39.264		
+	0.7836	44.775		
+	0.7837	50.423		
+	0.7838	56.289		
+	0.7839	62.217		
+	0.784	68.182		
+	0.7841	73.998		
+	0.7842	79.851		
+	0.7843	85.194		
+	0.7844	89.686		
+	0.7845	93.25		
+	0.7846	95.949		
+	0.7847	97.865		
+	0.7848	99.339		
+	0.7849	100.503		
+	0.785	101.286		
+	0.7851	101.865		
+	0.7852	102.45		
+	0.7853	103.016		
+	0.7854	103.501		
+	0.7855	104.21		
+	0.7856	104.994		
+	0.7857	105.678		
+	0.7858	106.362		
+	0.7859	107.239		
+	0.786	107.905		
+	0.7861	108.57		
+	0.7862	109.242		
+	0.7863	109.709		
+	0.7864	110.125		
+	0.7865	110.511		
+	0.7866	110.853		
+	0.7867	111.083		
+	0.7868	111.357		
+	0.7869	111.525		
+	0.787	111.575		
+	0.7871	111.724		
+	0.7872	111.879		
+	0.7873	111.96		
+	0.7874	111.879		
+	0.7875	111.848		
+	0.7876	111.991		
+	0.7877	112.035		
+	0.7878	111.985		
+	0.7879	112.11		
+	0.788	112.228		
+	0.7881	112.215		
+	0.7882	112.483		
+	0.7883	112.676		
+	0.7884	112.918		
+	0.7885	113.068		
+	0.7886	113.273		
+	0.7887	113.385		
+	0.7888	113.267		
+	0.7889	113.304		
+	0.789	113.117		
+	0.7891	112.452		
+	0.7892	111.68		
+	0.7893	110.461		
+	0.7894	108.62		
+	0.7895	106.138		
+	0.7896	102.779		
+	0.7897	98.058		
+	0.7898	91.066		
+	0.7899	81.904		
+	0.79	74.166		
+	0.7901	67.666		
+	0.7902	61.632		
+	0.7903	56.052		
+	0.7904	50.803		
+	0.7905	45.864		
+	0.7906	41.211		
+	0.7907	36.782		
+	0.7908	32.689		
+	0.7909	28.913		
+	0.791	25.331		
+	0.7911	21.86		
+	0.7912	18.681		
+	0.7913	15.789		
+	0.7914	13.052		
+	0.7915	10.557		
+	0.7916	8.343		
+	0.7917	6.346		
+	0.7918	4.567		
+	0.7919	2.981		
+	0.792	1.718		
+	0.7921	0.518		
+	0.7922	-0.378		
+	0.7923	-1.056		
+	0.7924	-1.765		
+	0.7925	-2.2		
+	0.7926	-2.505		
+	0.7927	-2.592		
+	0.7928	-2.847		
+	0.7929	-2.916		
+	0.793	-2.854		
+	0.7931	-2.841		
+	0.7932	-2.779		
+	0.7933	-2.667		
+	0.7934	-2.642		
+	0.7935	-2.555		
+	0.7936	-2.561		
+	0.7937	-2.356		
+	0.7938	-2.431		
+	0.7939	-2.381		
+	0.794	-2.238		
+	0.7941	-2.232		
+	0.7942	-2.281		
+	0.7943	-2.219		
+	0.7944	-2.113		
+	0.7945	-2.113		
+	0.7946	-2.101		
+	0.7947	-2.039		
+	0.7948	-1.989		
+	0.7949	-1.933		
+	0.795	-1.777		
+	0.7951	-1.759		
+	0.7952	-1.802		
+	0.7953	-1.634		
+	0.7954	-1.597		
+	0.7955	-1.622		
+	0.7956	-1.479		
+	0.7957	-1.491		
+	0.7958	-1.498		
+	0.7959	-1.473		
+	0.796	-1.448		
+	0.7961	-1.404		
+	0.7962	-1.361		
+	0.7963	-1.267		
+	0.7964	-1.062		
+	0.7965	-1.068		
+	0.7966	-0.938		
+	0.7967	-0.788		
+	0.7968	-0.708		
+	0.7969	-0.739		
+	0.797	-0.509		
+	0.7971	-0.49		
+	0.7972	-0.415		
+	0.7973	-0.278		
+	0.7974	-0.297		
+	0.7975	-0.322		
+	0.7976	-0.303		
+	0.7977	-0.222		
+	0.7978	-0.222		
+	0.7979	-0.235		
+	0.798	-0.179		
+	0.7981	-0.067		
+	0.7982	-0.216		
+	0.7983	0.039		
+	0.7984	0.219		
+	0.7985	0.344		
+	0.7986	0.717		
+	0.7987	1.382		
+	0.7988	2.222		
+	0.7989	3.678		
+	0.799	5.768		
+	0.7991	8.399		
+	0.7992	11.366		
+	0.7993	14.688		
+	0.7994	18.557		
+	0.7995	22.563		
+	0.7996	26.904		
+	0.7997	31.588		
+	0.7998	36.726		
+	0.7999	41.939		
+	0.8	47.636		
+	0.8001	53.421		
+	0.8002	59.212		
+	0.8003	65.184		
+	0.8004	71.249		
+	0.8005	76.99		
+	0.8006	82.576		
+	0.8007	87.533		
+	0.8008	91.595		
+	0.8009	94.568		
+	0.801	96.87		
+	0.8011	98.736		
+	0.8012	99.862		
+	0.8013	100.857		
+	0.8014	101.51		
+	0.8015	102.095		
+	0.8016	102.58		
+	0.8017	103.302		
+	0.8018	103.862		
+	0.8019	104.527		
+	0.802	105.386		
+	0.8021	106.2		
+	0.8022	106.872		
+	0.8023	107.693		
+	0.8024	108.396		
+	0.8025	108.968		
+	0.8026	109.454		
+	0.8027	110.076		
+	0.8028	110.393		
+	0.8029	110.635		
+	0.803	111.015		
+	0.8031	111.251		
+	0.8032	111.388		
+	0.8033	111.668		
+	0.8034	111.848		
+	0.8035	111.892		
+	0.8036	111.917		
+	0.8037	112.122		
+	0.8038	112.11		
+	0.8039	112.085		
+	0.804	112.24		
+	0.8041	112.215		
+	0.8042	112.153		
+	0.8043	112.203		
+	0.8044	112.402		
+	0.8045	112.514		
+	0.8046	112.607		
+	0.8047	112.837		
+	0.8048	113.074		
+	0.8049	113.18		
+	0.805	113.447		
+	0.8051	113.553		
+	0.8052	113.478		
+	0.8053	113.323		
+	0.8054	113.099		
+	0.8055	112.427		
+	0.8056	111.438		
+	0.8057	109.951		
+	0.8058	107.886		
+	0.8059	104.994		
+	0.806	101.199		
+	0.8061	95.993		
+	0.8062	87.508		
+	0.8063	78.701		
+	0.8064	71.703		
+	0.8065	65.433		
+	0.8066	59.443		
+	0.8067	54.186		
+	0.8068	49.117		
+	0.8069	44.147		
+	0.807	39.724		
+	0.8071	35.575		
+	0.8072	31.513		
+	0.8073	27.738		
+	0.8074	24.254		
+	0.8075	20.883		
+	0.8076	17.642		
+	0.8077	14.936		
+	0.8078	12.293		
+	0.8079	9.718		
+	0.808	7.609		
+	0.8081	5.755		
+	0.8082	3.951		
+	0.8083	2.477		
+	0.8084	1.407		
+	0.8085	0.281		
+	0.8086	-0.596		
+	0.8087	-1.143		
+	0.8088	-1.672		
+	0.8089	-2.207		
+	0.809	-2.406		
+	0.8091	-2.605		
+	0.8092	-2.816		
+	0.8093	-2.891		
+	0.8094	-2.754		
+	0.8095	-2.791		
+	0.8096	-2.866		
+	0.8097	-2.766		
+	0.8098	-2.611		
+	0.8099	-2.63		
+	0.81	-2.443		
+	0.8101	-2.35		
+	0.8102	-2.343		
+	0.8103	-2.269		
+	0.8104	-2.188		
+	0.8105	-2.138		
+	0.8106	-2.157		
+	0.8107	-2.088		
+	0.8108	-2.045		
+	0.8109	-2.057		
+	0.811	-2.07		
+	0.8111	-1.871		
+	0.8112	-1.914		
+	0.8113	-1.952		
+	0.8114	-1.79		
+	0.8115	-1.771		
+	0.8116	-1.883		
+	0.8117	-1.634		
+	0.8118	-1.498		
+	0.8119	-1.554		
+	0.812	-1.547		
+	0.8121	-1.33		
+	0.8122	-1.305		
+	0.8123	-1.342		
+	0.8124	-1.218		
+	0.8125	-1.211		
+	0.8126	-1.305		
+	0.8127	-1.068		
+	0.8128	-1.043		
+	0.8129	-1.012		
+	0.813	-0.956		
+	0.8131	-0.739		
+	0.8132	-0.67		
+	0.8133	-0.664		
+	0.8134	-0.397		
+	0.8135	-0.347		
+	0.8136	-0.39		
+	0.8137	-0.278		
+	0.8138	-0.104		
+	0.8139	-0.229		
+	0.814	-0.197		
+	0.8141	-0.067		
+	0.8142	-0.16		
+	0.8143	-0.26		
+	0.8144	-0.023		
+	0.8145	-0.017		
+	0.8146	-0.16		
+	0.8147	-0.104		
+	0.8148	0.25		
+	0.8149	0.418		
+	0.815	0.922		
+	0.8151	1.855		
+	0.8152	2.813		
+	0.8153	4.468		
+	0.8154	6.881		
+	0.8155	9.736		
+	0.8156	12.797		
+	0.8157	16.286		
+	0.8158	20.28		
+	0.8159	24.366		
+	0.816	28.764		
+	0.8161	33.678		
+	0.8162	38.692		
+	0.8163	44.035		
+	0.8164	49.801		
+	0.8165	55.648		
+	0.8166	61.433		
+	0.8167	67.479		
+	0.8168	73.463		
+	0.8169	79.08		
+	0.817	84.46		
+	0.8171	89.275		
+	0.8172	92.945		
+	0.8173	95.576		
+	0.8174	97.766		
+	0.8175	99.296		
+	0.8176	100.285		
+	0.8177	101.174		
+	0.8178	101.933		
+	0.8179	102.294		
+	0.818	102.736		
+	0.8181	103.526		
+	0.8182	104.123		
+	0.8183	104.77		
+	0.8184	105.703		
+	0.8185	106.53		
+	0.8186	107.177		
+	0.8187	108.004		
+	0.8188	108.701		
+	0.8189	109.261		
+	0.819	109.709		
+	0.8191	110.3		
+	0.8192	110.673		
+	0.8193	110.853		
+	0.8194	111.27		
+	0.8195	111.525		
+	0.8196	111.587		
+	0.8197	111.68		
+	0.8198	111.929		
+	0.8199	111.948		
+	0.82	112.06		
+	0.8201	112.228		
+	0.8202	112.253		
+	0.8203	112.166		
+	0.8204	112.321		
+	0.8205	112.495		
+	0.8206	112.464		
+	0.8207	112.508		
+	0.8208	112.682		
+	0.8209	112.738		
+	0.821	112.844		
+	0.8211	113.148		
+	0.8212	113.304		
+	0.8213	113.397		
+	0.8214	113.559		
+	0.8215	113.658		
+	0.8216	113.571		
+	0.8217	113.484		
+	0.8218	113.105		
+	0.8219	112.377		
+	0.822	111.22		
+	0.8221	109.715		
+	0.8222	107.569		
+	0.8223	104.403		
+	0.8224	100.235		
+	0.8225	94.369		
+	0.8226	85.257		
+	0.8227	76.94		
+	0.8228	70.291		
+	0.8229	64.021		
+	0.823	58.18		
+	0.8231	53.017		
+	0.8232	48.016		
+	0.8233	43.27		
+	0.8234	38.841		
+	0.8235	34.854		
+	0.8236	30.798		
+	0.8237	27.141		
+	0.8238	23.701		
+	0.8239	20.392		
+	0.824	17.226		
+	0.8241	14.476		
+	0.8242	11.92		
+	0.8243	9.369		
+	0.8244	7.236		
+	0.8245	5.444		
+	0.8246	3.659		
+	0.8247	2.179		
+	0.8248	1.115		
+	0.8249	0.132		
+	0.825	-0.764		
+	0.8251	-1.28		
+	0.8252	-1.777		
+	0.8253	-2.194		
+	0.8254	-2.431		
+	0.8255	-2.487		
+	0.8256	-2.729		
+	0.8257	-2.791		
+	0.8258	-2.717		
+	0.8259	-2.71		
+	0.826	-2.785		
+	0.8261	-2.661		
+	0.8262	-2.599		
+	0.8263	-2.623		
+	0.8264	-2.574		
+	0.8265	-2.424		
+	0.8266	-2.35		
+	0.8267	-2.256		
+	0.8268	-2.151		
+	0.8269	-2.138		
+	0.827	-2.12		
+	0.8271	-2.026		
+	0.8272	-1.945		
+	0.8273	-1.921		
+	0.8274	-1.889		
+	0.8275	-1.809		
+	0.8276	-1.939		
+	0.8277	-1.933		
+	0.8278	-1.771		
+	0.8279	-1.74		
+	0.828	-1.858		
+	0.8281	-1.697		
+	0.8282	-1.591		
+	0.8283	-1.56		
+	0.8284	-1.522		
+	0.8285	-1.274		
+	0.8286	-1.386		
+	0.8287	-1.305		
+	0.8288	-1.243		
+	0.8289	-1.149		
+	0.829	-1.174		
+	0.8291	-0.95		
+	0.8292	-0.963		
+	0.8293	-0.95		
+	0.8294	-0.863		
+	0.8295	-0.689		
+	0.8296	-0.645		
+	0.8297	-0.652		
+	0.8298	-0.502		
+	0.8299	-0.39		
+	0.83	-0.359		
+	0.8301	-0.247		
+	0.8302	-0.117		
+	0.8303	-0.104		
+	0.8304	-0.03		
+	0.8305	0.014		
+	0.8306	0.039		
+	0.8307	-0.054		
+	0.8308	0.026		
+	0.8309	-0.005		
+	0.831	-0.086		
+	0.8311	0.132		
+	0.8312	0.257		
+	0.8313	0.592		
+	0.8314	1.152		
+	0.8315	2.098		
+	0.8316	3.367		
+	0.8317	5.283		
+	0.8318	8.075		
+	0.8319	10.937		
+	0.832	14.19		
+	0.8321	17.891		
+	0.8322	21.99		
+	0.8323	26.164		
+	0.8324	30.755		
+	0.8325	35.675		
+	0.8326	40.769		
+	0.8327	46.243		
+	0.8328	51.904		
+	0.8329	57.763		
+	0.833	63.591		
+	0.8331	69.513		
+	0.8332	75.478		
+	0.8333	81.046		
+	0.8334	86.159		
+	0.8335	90.706		
+	0.8336	93.922		
+	0.8337	96.447		
+	0.8338	98.357		
+	0.8339	99.843		
+	0.834	100.727		
+	0.8341	101.448		
+	0.8342	102.145		
+	0.8343	102.524		
+	0.8344	103.04		
+	0.8345	103.718		
+	0.8346	104.266		
+	0.8347	104.875		
+	0.8348	105.84		
+	0.8349	106.717		
+	0.835	107.432		
+	0.8351	108.154		
+	0.8352	108.863		
+	0.8353	109.429		
+	0.8354	109.933		
+	0.8355	110.455		
+	0.8356	110.872		
+	0.8357	111.04		
+	0.8358	111.313		
+	0.8359	111.568		
+	0.836	111.68		
+	0.8361	111.799		
+	0.8362	111.96		
+	0.8363	111.998		
+	0.8364	112.035		
+	0.8365	112.153		
+	0.8366	112.246		
+	0.8367	112.321		
+	0.8368	112.483		
+	0.8369	112.502		
+	0.837	112.551		
+	0.8371	112.638		
+	0.8372	112.893		
+	0.8373	112.962		
+	0.8374	113.024		
+	0.8375	113.248		
+	0.8376	113.441		
+	0.8377	113.522		
+	0.8378	113.658		
+	0.8379	113.683		
+	0.838	113.503		
+	0.8381	113.242		
+	0.8382	112.912		
+	0.8383	112.166		
+	0.8384	110.872		
+	0.8385	109.248		
+	0.8386	106.773		
+	0.8387	103.463		
+	0.8388	98.966		
+	0.8389	92.242		
+	0.839	83.036		
+	0.8391	75.161		
+	0.8392	68.729		
+	0.8393	62.69		
+	0.8394	56.992		
+	0.8395	51.754		
+	0.8396	46.896		
+	0.8397	42.138		
+	0.8398	37.808		
+	0.8399	33.883		
+	0.84	29.977		
+	0.8401	26.382		
+	0.8402	22.936		
+	0.8403	19.776		
+	0.8404	16.728		
+	0.8405	13.991		
+	0.8406	11.459		
+	0.8407	9.033		
+	0.8408	6.9		
+	0.8409	5.065		
+	0.841	3.416		
+	0.8411	1.998		
+	0.8412	0.816		
+	0.8413	-0.092		
+	0.8414	-0.931		
+	0.8415	-1.479		
+	0.8416	-1.871		
+	0.8417	-2.269		
+	0.8418	-2.468		
+	0.8419	-2.549		
+	0.842	-2.648		
+	0.8421	-2.692		
+	0.8422	-2.592		
+	0.8423	-2.667		
+	0.8424	-2.667		
+	0.8425	-2.692		
+	0.8426	-2.567		
+	0.8427	-2.468		
+	0.8428	-2.505		
+	0.8429	-2.462		
+	0.843	-2.418		
+	0.8431	-2.381		
+	0.8432	-2.244		
+	0.8433	-2.12		
+	0.8434	-2.07		
+	0.8435	-2.039		
+	0.8436	-1.939		
+	0.8437	-1.877		
+	0.8438	-1.939		
+	0.8439	-1.777		
+	0.844	-1.815		
+	0.8441	-1.802		
+	0.8442	-1.79		
+	0.8443	-1.777		
+	0.8444	-1.703		
+	0.8445	-1.728		
+	0.8446	-1.641		
+	0.8447	-1.634		
+	0.8448	-1.628		
+	0.8449	-1.392		
+	0.845	-1.305		
+	0.8451	-1.249		
+	0.8452	-1.28		
+	0.8453	-1.05		
+	0.8454	-0.987		
+	0.8455	-0.907		
+	0.8456	-0.851		
+	0.8457	-0.826		
+	0.8458	-0.832		
+	0.8459	-0.683		
+	0.846	-0.633		
+	0.8461	-0.533		
+	0.8462	-0.459		
+	0.8463	-0.378		
+	0.8464	-0.309		
+	0.8465	-0.291		
+	0.8466	-0.092		
+	0.8467	-0.117		
+	0.8468	-0.042		
+	0.8469	0.026		
+	0.847	0.07		
+	0.8471	0.051		
+	0.8472	0.138		
+	0.8473	0.12		
+	0.8474	0.145		
+	0.8475	0.163		
+	0.8476	0.437		
+	0.8477	0.866		
+	0.8478	1.414		
+	0.8479	2.371		
+	0.848	3.908		
+	0.8481	6.085		
+	0.8482	8.853		
+	0.8483	11.969		
+	0.8484	15.316		
+	0.8485	19.166		
+	0.8486	23.253		
+	0.8487	27.607		
+	0.8488	32.235		
+	0.8489	37.255		
+	0.849	42.474		
+	0.8491	47.96		
+	0.8492	53.651		
+	0.8493	59.48		
+	0.8494	65.358		
+	0.8495	71.093		
+	0.8496	76.89		
+	0.8497	82.439		
+	0.8498	87.365		
+	0.8499	91.527		
+	0.85	94.668		
+	0.8501	96.988		
+	0.8502	98.674		
+	0.8503	100.061		
+	0.8504	100.95		
+	0.8505	101.604		
+	0.8506	102.232		
+	0.8507	102.773		
+	0.8508	103.24		
+	0.8509	103.762		
+	0.851	104.465		
+	0.8511	105.168		
+	0.8512	105.871		
+	0.8513	106.779		
+	0.8514	107.5		
+	0.8515	108.203		
+	0.8516	108.863		
+	0.8517	109.534		
+	0.8518	110.038		
+	0.8519	110.443		
+	0.852	110.785		
+	0.8521	111.108		
+	0.8522	111.425		
+	0.8523	111.618		
+	0.8524	111.799		
+	0.8525	111.861		
+	0.8526	111.917		
+	0.8527	112.097		
+	0.8528	112.035		
+	0.8529	112.041		
+	0.853	112.172		
+	0.8531	112.24		
+	0.8532	112.315		
+	0.8533	112.446		
+	0.8534	112.595		
+	0.8535	112.669		
+	0.8536	112.806		
+	0.8537	112.999		
+	0.8538	113.155		
+	0.8539	113.291		
+	0.854	113.59		
+	0.8541	113.652		
+	0.8542	113.584		
+	0.8543	113.683		
+	0.8544	113.615		
+	0.8545	113.192		
+	0.8546	112.669		
+	0.8547	111.805		
+	0.8548	110.461		
+	0.8549	108.57		
+	0.855	106.132		
+	0.8551	102.63		
+	0.8552	97.66		
+	0.8553	90.227		
+	0.8554	81.307		
+	0.8555	73.886		
+	0.8556	67.467		
+	0.8557	61.576		
+	0.8558	55.978		
+	0.8559	50.803		
+	0.856	45.976		
+	0.8561	41.422		
+	0.8562	37.062		
+	0.8563	33.093		
+	0.8564	29.305		
+	0.8565	25.704		
+	0.8566	22.382		
+	0.8567	19.26		
+	0.8568	16.212		
+	0.8569	13.5		
+	0.857	11.036		
+	0.8571	8.753		
+	0.8572	6.744		
+	0.8573	4.853		
+	0.8574	3.329		
+	0.8575	1.855		
+	0.8576	0.661		
+	0.8577	-0.142		
+	0.8578	-1.019		
+	0.8579	-1.609		
+	0.858	-1.976		
+	0.8581	-2.275		
+	0.8582	-2.561		
+	0.8583	-2.592		
+	0.8584	-2.636		
+	0.8585	-2.661		
+	0.8586	-2.679		
+	0.8587	-2.555		
+	0.8588	-2.543		
+	0.8589	-2.58		
+	0.859	-2.468		
+	0.8591	-2.462		
+	0.8592	-2.53		
+	0.8593	-2.431		
+	0.8594	-2.281		
+	0.8595	-2.343		
+	0.8596	-2.288		
+	0.8597	-2.207		
+	0.8598	-2.144		
+	0.8599	-2.07		
+	0.86	-1.964		
+	0.8601	-1.827		
+	0.8602	-1.908		
+	0.8603	-1.802		
+	0.8604	-1.634		
+	0.8605	-1.684		
+	0.8606	-1.728		
+	0.8607	-1.634		
+	0.8608	-1.684		
+	0.8609	-1.703		
+	0.861	-1.609		
+	0.8611	-1.485		
+	0.8612	-1.541		
+	0.8613	-1.485		
+	0.8614	-1.354		
+	0.8615	-1.342		
+	0.8616	-1.267		
+	0.8617	-1.019		
+	0.8618	-0.95		
+	0.8619	-0.981		
+	0.862	-0.857		
+	0.8621	-0.658		
+	0.8622	-0.633		
+	0.8623	-0.614		
+	0.8624	-0.477		
+	0.8625	-0.49		
+	0.8626	-0.502		
+	0.8627	-0.285		
+	0.8628	-0.229		
+	0.8629	-0.297		
+	0.863	-0.117		
+	0.8631	-0.061		
+	0.8632	-0.079		
+	0.8633	0.014		
+	0.8634	0.176		
+	0.8635	0.107		
+	0.8636	0.002		
+	0.8637	0.244		
+	0.8638	0.275		
+	0.8639	0.294		
+	0.864	0.586		
+	0.8641	1.078		
+	0.8642	1.582		
+	0.8643	2.608		
+	0.8644	4.231		
+	0.8645	6.489		
+	0.8646	9.145		
+	0.8647	12.311		
+	0.8648	15.751		
+	0.8649	19.533		
+	0.865	23.726		
+	0.8651	28.204		
+	0.8652	32.789		
+	0.8653	37.821		
+	0.8654	43.22		
+	0.8655	48.719		
+	0.8656	54.261		
+	0.8657	60.158		
+	0.8658	65.968		
+	0.8659	71.709		
+	0.866	77.432		
+	0.8661	83.024		
+	0.8662	87.745		
+	0.8663	91.614		
+	0.8664	94.73		
+	0.8665	96.963		
+	0.8666	98.637		
+	0.8667	100.024		
+	0.8668	100.957		
+	0.8669	101.529		
+	0.867	102.139		
+	0.8671	102.736		
+	0.8672	103.296		
+	0.8673	103.756		
+	0.8674	104.564		
+	0.8675	105.168		
+	0.8676	105.858		
+	0.8677	106.773		
+	0.8678	107.55		
+	0.8679	108.079		
+	0.868	108.763		
+	0.8681	109.354		
+	0.8682	109.845		
+	0.8683	110.206		
+	0.8684	110.704		
+	0.8685	111.034		
+	0.8686	111.208		
+	0.8687	111.568		
+	0.8688	111.805		
+	0.8689	111.855		
+	0.869	111.979		
+	0.8691	112.06		
+	0.8692	112.004		
+	0.8693	112.016		
+	0.8694	112.209		
+	0.8695	112.166		
+	0.8696	112.135		
+	0.8697	112.253		
+	0.8698	112.458		
+	0.8699	112.446		
+	0.87	112.657		
+	0.8701	112.949		
+	0.8702	113.03		
+	0.8703	113.211		
+	0.8704	113.478		
+	0.8705	113.646		
+	0.8706	113.615		
+	0.8707	113.652		
+	0.8708	113.503		
+	0.8709	113.148		
+	0.871	112.427		
+	0.8711	111.73		
+	0.8712	110.188		
+	0.8713	108.253		
+	0.8714	105.703		
+	0.8715	102.257		
+	0.8716	97.262		
+	0.8717	89.654		
+	0.8718	80.934		
+	0.8719	73.42		
+	0.872	67.143		
+	0.8721	61.445		
+	0.8722	55.853		
+	0.8723	50.647		
+	0.8724	45.864		
+	0.8725	41.248		
+	0.8726	36.844		
+	0.8727	32.975		
+	0.8728	29.231		
+	0.8729	25.449		
+	0.873	22.121		
+	0.8731	19.129		
+	0.8732	16.143		
+	0.8733	13.369		
+	0.8734	10.949		
+	0.8735	8.797		
+	0.8736	6.614		
+	0.8737	4.835		
+	0.8738	3.348		
+	0.8739	1.899		
+	0.874	0.785		
+	0.8741	-0.148		
+	0.8742	-0.944		
+	0.8743	-1.597		
+	0.8744	-1.927		
+	0.8745	-2.244		
+	0.8746	-2.679		
+	0.8747	-2.686		
+	0.8748	-2.661		
+	0.8749	-2.717		
+	0.875	-2.723		
+	0.8751	-2.549		
+	0.8752	-2.561		
+	0.8753	-2.605		
+	0.8754	-2.462		
+	0.8755	-2.337		
+	0.8756	-2.424		
+	0.8757	-2.325		
+	0.8758	-2.194		
+	0.8759	-2.238		
+	0.876	-2.281		
+	0.8761	-2.095		
+	0.8762	-2.151		
+	0.8763	-2.169		
+	0.8764	-1.995		
+	0.8765	-1.889		
+	0.8766	-1.896		
+	0.8767	-1.858		
+	0.8768	-1.616		
+	0.8769	-1.672		
+	0.877	-1.659		
+	0.8771	-1.498		
+	0.8772	-1.466		
+	0.8773	-1.609		
+	0.8774	-1.491		
+	0.8775	-1.41		
+	0.8776	-1.516		
+	0.8777	-1.485		
+	0.8778	-1.261		
+	0.8779	-1.354		
+	0.878	-1.305		
+	0.8781	-1.093		
+	0.8782	-0.95		
+	0.8783	-0.907		
+	0.8784	-0.77		
+	0.8785	-0.558		
+	0.8786	-0.583		
+	0.8787	-0.564		
+	0.8788	-0.359		
+	0.8789	-0.316		
+	0.879	-0.39		
+	0.8791	-0.272		
+	0.8792	-0.185		
+	0.8793	-0.26		
+	0.8794	-0.098		
+	0.8795	0.014		
+	0.8796	-0.086		
+	0.8797	-0.086		
+	0.8798	0.114		
+	0.8799	0.107		
+	0.88	0.002		
+	0.8801	0.294		
+	0.8802	0.294		
+	0.8803	0.319		
+	0.8804	0.692		
+	0.8805	1.264		
+	0.8806	1.855		
+	0.8807	2.906		
+	0.8808	4.692		
+	0.8809	7.074		
+	0.881	9.693		
+	0.8811	12.996		
+	0.8812	16.454		
+	0.8813	20.224		
+	0.8814	24.447		
+	0.8815	28.951		
+	0.8816	33.566		
+	0.8817	38.611		
+	0.8818	44.122		
+	0.8819	49.583		
+	0.882	55.194		
+	0.8821	61.066		
+	0.8822	66.963		
+	0.8823	72.574		
+	0.8824	78.284		
+	0.8825	83.615		
+	0.8826	88.218		
+	0.8827	91.9		
+	0.8828	94.898		
+	0.8829	96.976		
+	0.883	98.5		
+	0.8831	99.793		
+	0.8832	100.739		
+	0.8833	101.305		
+	0.8834	101.971		
+	0.8835	102.605		
+	0.8836	103.022		
+	0.8837	103.712		
+	0.8838	104.484		
+	0.8839	105.205		
+	0.884	105.877		
+	0.8841	106.704		
+	0.8842	107.401		
+	0.8843	107.948		
+	0.8844	108.601		
+	0.8845	109.286		
+	0.8846	109.653		
+	0.8847	109.933		
+	0.8848	110.436		
+	0.8849	110.754		
+	0.885	110.996		
+	0.8851	111.351		
+	0.8852	111.581		
+	0.8853	111.6		
+	0.8854	111.761		
+	0.8855	111.929		
+	0.8856	111.867		
+	0.8857	111.848		
+	0.8858	111.935		
+	0.8859	112.004		
+	0.886	111.917		
+	0.8861	112.066		
+	0.8862	112.178		
+	0.8863	112.215		
+	0.8864	112.296		
+	0.8865	112.607		
+	0.8866	112.806		
+	0.8867	112.937		
+	0.8868	113.279		
+	0.8869	113.366		
+	0.887	113.291		
+	0.8871	113.397		
+	0.8872	113.229		
+	0.8873	112.781		
+	0.8874	112.122		
+	0.8875	111.201		
+	0.8876	109.696		
+	0.8877	107.606		
+	0.8878	104.907		
+	0.8879	101.162		
+	0.888	95.9		
+	0.8881	87.813		
+	0.8882	79.291		
+	0.8883	72.132		
+	0.8884	66.017		
+	0.8885	60.326		
+	0.8886	54.889		
+	0.8887	49.776		
+	0.8888	44.993		
+	0.8889	40.452		
+	0.889	36.197		
+	0.8891	32.279		
+	0.8892	28.584		
+	0.8893	24.97		
+	0.8894	21.567		
+	0.8895	18.538		
+	0.8896	15.633		
+	0.8897	12.772		
+	0.8898	10.483		
+	0.8899	8.349		
+	0.89	6.259		
+	0.8901	4.586		
+	0.8902	3.056		
+	0.8903	1.725		
+	0.8904	0.636		
+	0.8905	-0.229		
+	0.8906	-0.95		
+	0.8907	-1.634		
+	0.8908	-2.07		
+	0.8909	-2.312		
+	0.891	-2.605		
+	0.8911	-2.698		
+	0.8912	-2.71		
+	0.8913	-2.76		
+	0.8914	-2.829		
+	0.8915	-2.636		
+	0.8916	-2.617		
+	0.8917	-2.549		
+	0.8918	-2.381		
+	0.8919	-2.368		
+	0.892	-2.387		
+	0.8921	-2.312		
+	0.8922	-2.213		
+	0.8923	-2.176		
+	0.8924	-2.219		
+	0.8925	-2.132		
+	0.8926	-2.088		
+	0.8927	-2.132		
+	0.8928	-2.02		
+	0.8929	-1.933		
+	0.893	-1.939		
+	0.8931	-1.889		
+	0.8932	-1.734		
+	0.8933	-1.728		
+	0.8934	-1.684		
+	0.8935	-1.535		
+	0.8936	-1.522		
+	0.8937	-1.491		
+	0.8938	-1.41		
+	0.8939	-1.379		
+	0.894	-1.435		
+	0.8941	-1.41		
+	0.8942	-1.323		
+	0.8943	-1.354		
+	0.8944	-1.236		
+	0.8945	-1.124		
+	0.8946	-0.987		
+	0.8947	-1.006		
+	0.8948	-0.888		
+	0.8949	-0.708		
+	0.895	-0.664		
+	0.8951	-0.54		
+	0.8952	-0.428		
+	0.8953	-0.347		
+	0.8954	-0.341		
+	0.8955	-0.197		
+	0.8956	-0.061		
+	0.8957	-0.098		
+	0.8958	-0.11		
+	0.8959	0.008		
+	0.896	-0.005		
+	0.8961	-0.023		
+	0.8962	0.045		
+	0.8963	0.089		
+	0.8964	-0.048		
+	0.8965	0.138		
+	0.8966	0.194		
+	0.8967	0.362		
+	0.8968	0.686		
+	0.8969	1.183		
+	0.897	1.917		
+	0.8971	3.006		
+	0.8972	4.853		
+	0.8973	7.205		
+	0.8974	9.91		
+	0.8975	13.014		
+	0.8976	16.597		
+	0.8977	20.448		
+	0.8978	24.547		
+	0.8979	29.038		
+	0.898	33.722		
+	0.8981	38.679		
+	0.8982	44.141		
+	0.8983	49.614		
+	0.8984	55.331		
+	0.8985	61.134		
+	0.8986	66.919		
+	0.8987	72.654		
+	0.8988	78.284		
+	0.8989	83.639		
+	0.899	88.224		
+	0.8991	91.819		
+	0.8992	94.649		
+	0.8993	96.808		
+	0.8994	98.413		
+	0.8995	99.563		
+	0.8996	100.459		
+	0.8997	101.125		
+	0.8998	101.647		
+	0.8999	102.275		
+	0.9	102.81		
+	0.9001	103.501		
+	0.9002	104.191		
+	0.9003	104.987		
+	0.9004	105.74		
+	0.9005	106.499		
+	0.9006	107.295		
+	0.9007	107.892		
+	0.9008	108.415		
+	0.9009	109.018		
+	0.901	109.472		
+	0.9011	109.833		
+	0.9012	110.138		
+	0.9013	110.486		
+	0.9014	110.735		
+	0.9015	110.978		
+	0.9016	111.251		
+	0.9017	111.425		
+	0.9018	111.6		
+	0.9019	111.674		
+	0.902	111.73		
+	0.9021	111.68		
+	0.9022	111.811		
+	0.9023	111.83		
+	0.9024	111.811		
+	0.9025	111.861		
+	0.9026	111.973		
+	0.9027	112.116		
+	0.9028	112.147		
+	0.9029	112.352		
+	0.903	112.564		
+	0.9031	112.669		
+	0.9032	112.974		
+	0.9033	113.117		
+	0.9034	113.148		
+	0.9035	113.167		
+	0.9036	113.049		
+	0.9037	112.638		
+	0.9038	111.935		
+	0.9039	111.046		
+	0.904	109.584		
+	0.9041	107.413		
+	0.9042	104.714		
+	0.9043	100.988		
+	0.9044	95.763		
+	0.9045	87.633		
+	0.9046	79.018		
+	0.9047	72.014		
+	0.9048	65.762		
+	0.9049	60.065		
+	0.905	54.703		
+	0.9051	49.72		
+	0.9052	44.868		
+	0.9053	40.458		
+	0.9054	36.21		
+	0.9055	32.291		
+	0.9056	28.596		
+	0.9057	25.032		
+	0.9058	21.648		
+	0.9059	18.47		
+	0.906	15.633		
+	0.9061	12.846		
+	0.9062	10.402		
+	0.9063	8.256		
+	0.9064	6.216		
+	0.9065	4.499		
+	0.9066	3.012		
+	0.9067	1.774		
+	0.9068	0.617		
+	0.9069	-0.247		
+	0.907	-0.925		
+	0.9071	-1.535		
+	0.9072	-2.001		
+	0.9073	-2.238		
+	0.9074	-2.48		
+	0.9075	-2.617		
+	0.9076	-2.704		
+	0.9077	-2.673		
+	0.9078	-2.735		
+	0.9079	-2.729		
+	0.908	-2.642		
+	0.9081	-2.648		
+	0.9082	-2.58		
+	0.9083	-2.387		
+	0.9084	-2.406		
+	0.9085	-2.294		
+	0.9086	-2.219		
+	0.9087	-2.151		
+	0.9088	-2.088		
+	0.9089	-2.057		
+	0.909	-2.02		
+	0.9091	-2.045		
+	0.9092	-2.057		
+	0.9093	-1.958		
+	0.9094	-1.871		
+	0.9095	-1.871		
+	0.9096	-1.833		
+	0.9097	-1.765		
+	0.9098	-1.721		
+	0.9099	-1.697		
+	0.91	-1.572		
+	0.9101	-1.473		
+	0.9102	-1.491		
+	0.9103	-1.348		
+	0.9104	-1.373		
+	0.9105	-1.336		
+	0.9106	-1.274		
+	0.9107	-1.174		
+	0.9108	-1.18		
+	0.9109	-1.124		
+	0.911	-1.006		
+	0.9111	-0.931		
+	0.9112	-0.931		
+	0.9113	-0.764		
+	0.9114	-0.714		
+	0.9115	-0.664		
+	0.9116	-0.453		
+	0.9117	-0.322		
+	0.9118	-0.229		
+	0.9119	-0.191		
+	0.912	-0.086		
+	0.9121	0.045		
+	0.9122	-0.042		
+	0.9123	0.082		
+	0.9124	0.051		
+	0.9125	-0.005		
+	0.9126	0.002		
+	0.9127	0.114		
+	0.9128	0.008		
+	0.9129	0.008		
+	0.913	0.163		
+	0.9131	0.331		
+	0.9132	0.648		
+	0.9133	1.227		
+	0.9134	2.104		
+	0.9135	3.23		
+	0.9136	5.127		
+	0.9137	7.628		
+	0.9138	10.433		
+	0.9139	13.668		
+	0.914	17.201		
+	0.9141	21.076		
+	0.9142	25.088		
+	0.9143	29.56		
+	0.9144	34.437		
+	0.9145	39.376		
+	0.9146	44.638		
+	0.9147	50.23		
+	0.9148	55.897		
+	0.9149	61.545		
+	0.915	67.442		
+	0.9151	73.214		
+	0.9152	78.676		
+	0.9153	83.975		
+	0.9154	88.504		
+	0.9155	92.043		
+	0.9156	94.78		
+	0.9157	96.907		
+	0.9158	98.406		
+	0.9159	99.538		
+	0.916	100.378		
+	0.9161	101.137		
+	0.9162	101.548		
+	0.9163	102.157		
+	0.9164	102.748		
+	0.9165	103.364		
+	0.9166	104.048		
+	0.9167	104.931		
+	0.9168	105.709		
+	0.9169	106.399		
+	0.917	107.227		
+	0.9171	107.923		
+	0.9172	108.421		
+	0.9173	108.993		
+	0.9174	109.466		
+	0.9175	109.733		
+	0.9176	109.989		
+	0.9177	110.43		
+	0.9178	110.673		
+	0.9179	110.797		
+	0.918	111.065		
+	0.9181	111.245		
+	0.9182	111.394		
+	0.9183	111.481		
+	0.9184	111.668		
+	0.9185	111.6		
+	0.9186	111.568		
+	0.9187	111.755		
+	0.9188	111.792		
+	0.9189	111.799		
+	0.919	111.973		
+	0.9191	112.091		
+	0.9192	112.023		
+	0.9193	112.203		
+	0.9194	112.489		
+	0.9195	112.576		
+	0.9196	112.707		
+	0.9197	112.962		
+	0.9198	112.931		
+	0.9199	112.875		
+	0.92	112.781		
+	0.9201	112.446		
+	0.9202	111.705		
+	0.9203	110.704		
+	0.9204	109.217		
+	0.9205	107.077		
+	0.9206	104.185		
+	0.9207	100.403		
+	0.9208	94.911		
+	0.9209	86.364		
+	0.921	78.029		
+	0.9211	71.255		
+	0.9212	64.979		
+	0.9213	59.281		
+	0.9214	54.087		
+	0.9215	49.055		
+	0.9216	44.277		
+	0.9217	40.004		
+	0.9218	35.874		
+	0.9219	31.806		
+	0.922	28.155		
+	0.9221	24.74		
+	0.9222	21.368		
+	0.9223	18.19		
+	0.9224	15.484		
+	0.9225	12.678		
+	0.9226	10.11		
+	0.9227	8.051		
+	0.9228	6.06		
+	0.9229	4.275		
+	0.923	2.788		
+	0.9231	1.55		
+	0.9232	0.449		
+	0.9233	-0.453		
+	0.9234	-0.938		
+	0.9235	-1.541		
+	0.9236	-2.039		
+	0.9237	-2.263		
+	0.9238	-2.437		
+	0.9239	-2.636		
+	0.924	-2.648		
+	0.9241	-2.692		
+	0.9242	-2.71		
+	0.9243	-2.798		
+	0.9244	-2.605		
+	0.9245	-2.599		
+	0.9246	-2.623		
+	0.9247	-2.518		
+	0.9248	-2.412		
+	0.9249	-2.387		
+	0.925	-2.238		
+	0.9251	-2.132		
+	0.9252	-2.157		
+	0.9253	-2.132		
+	0.9254	-2.001		
+	0.9255	-1.889		
+	0.9256	-1.983		
+	0.9257	-1.877		
+	0.9258	-1.827		
+	0.9259	-1.908		
+	0.926	-1.833		
+	0.9261	-1.74		
+	0.9262	-1.79		
+	0.9263	-1.815		
+	0.9264	-1.684		
+	0.9265	-1.529		
+	0.9266	-1.616		
+	0.9267	-1.386		
+	0.9268	-1.286		
+	0.9269	-1.429		
+	0.927	-1.286		
+	0.9271	-1.099		
+	0.9272	-1.081		
+	0.9273	-0.994		
+	0.9274	-0.963		
+	0.9275	-0.894		
+	0.9276	-0.931		
+	0.9277	-0.795		
+	0.9278	-0.652		
+	0.9279	-0.658		
+	0.928	-0.614		
+	0.9281	-0.384		
+	0.9282	-0.316		
+	0.9283	-0.297		
+	0.9284	-0.017		
+	0.9285	0.064		
+	0.9286	-0.036		
+	0.9287	0.12		
+	0.9288	0.201		
+	0.9289	0.051		
+	0.929	0.089		
+	0.9291	0.145		
+	0.9292	0.17		
+	0.9293	0.014		
+	0.9294	0.188		
+	0.9295	0.431		
+	0.9296	0.58		
+	0.9297	1.14		
+	0.9298	1.98		
+	0.9299	3.112		
+	0.93	4.878		
+	0.9301	7.509		
+	0.9302	10.178		
+	0.9303	13.245		
+	0.9304	16.89		
+	0.9305	20.715		
+	0.9306	24.802		
+	0.9307	29.2		
+	0.9308	33.946		
+	0.9309	38.86		
+	0.931	44.047		
+	0.9311	49.664		
+	0.9312	55.163		
+	0.9313	60.836		
+	0.9314	66.733		
+	0.9315	72.381		
+	0.9316	77.917		
+	0.9317	83.254		
+	0.9318	87.975		
+	0.9319	91.508		
+	0.932	94.326		
+	0.9321	96.59		
+	0.9322	98.151		
+	0.9323	99.252		
+	0.9324	100.248		
+	0.9325	100.95		
+	0.9326	101.386		
+	0.9327	101.971		
+	0.9328	102.605		
+	0.9329	103.103		
+	0.933	103.768		
+	0.9331	104.62		
+	0.9332	105.441		
+	0.9333	106.107		
+	0.9334	107.009		
+	0.9335	107.724		
+	0.9336	108.234		
+	0.9337	108.8		
+	0.9338	109.36		
+	0.9339	109.715		
+	0.934	109.989		
+	0.9341	110.318		
+	0.9342	110.573		
+	0.9343	110.66		
+	0.9344	110.99		
+	0.9345	111.201		
+	0.9346	111.226		
+	0.9347	111.307		
+	0.9348	111.5		
+	0.9349	111.544		
+	0.935	111.544		
+	0.9351	111.674		
+	0.9352	111.743		
+	0.9353	111.761		
+	0.9354	111.886		
+	0.9355	112.06		
+	0.9356	112.128		
+	0.9357	112.178		
+	0.9358	112.47		
+	0.9359	112.545		
+	0.936	112.57		
+	0.9361	112.9		
+	0.9362	112.887		
+	0.9363	112.819		
+	0.9364	112.663		
+	0.9365	112.458		
+	0.9366	111.73		
+	0.9367	110.772		
+	0.9368	109.441		
+	0.9369	107.395		
+	0.937	104.596		
+	0.9371	101.131		
+	0.9372	95.999		
+	0.9373	87.981		
+	0.9374	79.391		
+	0.9375	72.35		
+	0.9376	66.036		
+	0.9377	60.32		
+	0.9378	54.964		
+	0.9379	49.894		
+	0.938	45.092		
+	0.9381	40.645		
+	0.9382	36.533		
+	0.9383	32.459		
+	0.9384	28.851		
+	0.9385	25.436		
+	0.9386	22.04		
+	0.9387	18.868		
+	0.9388	16.031		
+	0.9389	13.288		
+	0.939	10.744		
+	0.9391	8.579		
+	0.9392	6.508		
+	0.9393	4.623		
+	0.9394	3.124		
+	0.9395	1.874		
+	0.9396	0.611		
+	0.9397	-0.316		
+	0.9398	-0.894		
+	0.9399	-1.498		
+	0.94	-2.026		
+	0.9401	-2.207		
+	0.9402	-2.387		
+	0.9403	-2.549		
+	0.9404	-2.599		
+	0.9405	-2.518		
+	0.9406	-2.648		
+	0.9407	-2.655		
+	0.9408	-2.518		
+	0.9409	-2.536		
+	0.941	-2.63		
+	0.9411	-2.48		
+	0.9412	-2.399		
+	0.9413	-2.449		
+	0.9414	-2.443		
+	0.9415	-2.151		
+	0.9416	-2.219		
+	0.9417	-2.12		
+	0.9418	-1.952		
+	0.9419	-1.983		
+	0.942	-1.958		
+	0.9421	-1.846		
+	0.9422	-1.746		
+	0.9423	-1.79		
+	0.9424	-1.796		
+	0.9425	-1.715		
+	0.9426	-1.784		
+	0.9427	-1.715		
+	0.9428	-1.672		
+	0.9429	-1.628		
+	0.943	-1.603		
+	0.9431	-1.504		
+	0.9432	-1.361		
+	0.9433	-1.404		
+	0.9434	-1.224		
+	0.9435	-1.087		
+	0.9436	-1.093		
+	0.9437	-1.019		
+	0.9438	-0.863		
+	0.9439	-0.813		
+	0.944	-0.776		
+	0.9441	-0.708		
+	0.9442	-0.558		
+	0.9443	-0.664		
+	0.9444	-0.527		
+	0.9445	-0.341		
+	0.9446	-0.372		
+	0.9447	-0.291		
+	0.9448	-0.148		
+	0.9449	-0.067		
+	0.945	0.008		
+	0.9451	0.101		
+	0.9452	0.157		
+	0.9453	0.157		
+	0.9454	0.176		
+	0.9455	0.306		
+	0.9456	0.225		
+	0.9457	0.176		
+	0.9458	0.294		
+	0.9459	0.418		
+	0.946	0.53		
+       r       0				
.ends				
